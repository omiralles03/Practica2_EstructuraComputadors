//: version "1.8.7"

module CONTROL(Jump, MemWrite, ALUOp, ALUSrc, RegWrite, MemRead, Branch, MemToReg, funct, op, RegDst);
//: interface  /sz:(148, 230) /bd:[ Li0>op[5:0](142/230) Li1>funct[5:0](187/230) Ro0<RegWrite(201/230) Ro1<ALUSrc(174/230) Ro2<ALUOp[3:0](137/230) Ro3<MemToReg(115/230) Ro4<MemRead(89/230) Ro5<Branch(66/230) Ro6<Jump(43/230) Ro7<RegDst(23/230) Ro8<MemWrite(158/230) ]
output Branch;    //: /sn:0 /dp:15 {0}(1075,393)(936,393){1}
//: {2}(934,391)(934,331){3}
//: {4}(936,329)(1023,329){5}
//: {6}(934,327)(934,285)(1023,285){7}
//: {8}(934,395)(934,476){9}
//: {10}(932,478)(923,478)(923,465){11}
//: {12}(934,480)(934,498)(446,498)(446,347){13}
//: {14}(448,345)(570,345){15}
//: {16}(446,343)(446,283){17}
//: {18}(446,279)(446,252){19}
//: {20}(444,281)(417,281)(417,273){21}
supply0 w3;    //: /sn:0 {0}(1150,376)(1129,376)(1129,393){1}
output MemWrite;    //: /sn:0 {0}(571,423)(380,423){1}
//: {2}(378,421)(378,285){3}
//: {4}(378,281)(378,254){5}
//: {6}(376,283)(362,283)(362,275){7}
//: {8}(378,425)(378,441)(525,441){9}
output ALUSrc;    //: /sn:0 {0}(571,444)(546,444){1}
output RegDst;    //: /sn:0 {0}(1023,334)(959,334){1}
//: {2}(957,332)(957,290)(1023,290){3}
//: {4}(957,336)(957,356){5}
//: {6}(959,358)(1071,358){7}
//: {8}(957,360)(957,410){9}
//: {10}(959,412)(1026,412){11}
//: {12}(957,414)(957,477){13}
//: {14}(959,479)(974,479)(974,471){15}
//: {16}(957,481)(957,514)(238,514)(238,472){17}
//: {18}(240,470)(524,470){19}
//: {20}(238,468)(238,296){21}
//: {22}(240,294)(570,294){23}
//: {24}(238,292)(238,252){25}
//: {26}(236,294)(215,294)(215,270){27}
output RegWrite;    //: /sn:0 /dp:1 {0}(545,468)(572,468){1}
output [3:0] ALUOp;    //: /sn:0 {0}(1156,361)(1168,361){1}
//: {2}(1172,361)(1191,361){3}
//: {4}(1170,363)(1170,392){5}
output MemRead;    //: /sn:0 /dp:1 {0}(307,103)(307,89)(334,89)(334,371)(570,371){1}
input [5:0] funct;    //: /sn:0 {0}(911,468)(898,468){1}
//: {2}(897,468)(880,468){3}
//: {4}(879,468)(860,468){5}
//: {6}(859,468)(840,468){7}
//: {8}(839,468)(826,468){9}
//: {10}(824,466)(824,417)(818,417){11}
//: {12}(822,468)(809,468){13}
output MemToReg;    //: /sn:0 /dp:1 {0}(570,392)(310,392){1}
//: {2}(308,390)(308,287){3}
//: {4}(308,283)(308,254){5}
//: {6}(306,285)(294,285)(294,274){7}
//: {8}(308,394)(308,444){9}
//: {10}(310,446)(525,446){11}
//: {12}(308,448)(308,465)(524,465){13}
input [5:0] op;    //: /sn:0 {0}(149,177)(185,177){1}
output Jump;    //: /sn:0 {0}(571,320)(507,320)(507,284){1}
//: {2}(507,280)(507,252){3}
//: {4}(505,282)(486,282)(486,274){5}
wire w6;    //: /sn:0 {0}(1092,319)(1113,319)(1113,346)(1150,346){1}
wire w7;    //: /sn:0 {0}(250,231)(250,204){1}
//: {2}(252,202)(318,202){3}
//: {4}(322,202)(388,202){5}
//: {6}(392,202)(456,202){7}
//: {8}(460,202)(517,202){9}
//: {10}(521,202)(665,202){11}
//: {12}(519,204)(519,231){13}
//: {14}(458,204)(458,231){15}
//: {16}(390,204)(390,233){17}
//: {18}(320,200)(320,124){19}
//: {20}(320,204)(320,233){21}
//: {22}(248,202)(191,202){23}
wire w4;    //: /sn:0 {0}(1092,356)(1150,356){1}
wire w39;    //: /sn:0 {0}(504,231)(504,174){1}
//: {2}(506,172)(665,172){3}
//: {4}(502,172)(445,172){5}
//: {6}(441,172)(377,172){7}
//: {8}(373,172)(307,172){9}
//: {10}(305,170)(305,124){11}
//: {12}(303,172)(237,172){13}
//: {14}(233,172)(191,172){15}
//: {16}(235,174)(235,231){17}
//: {18}(305,174)(305,233){19}
//: {20}(375,174)(375,233){21}
//: {22}(443,174)(443,231){23}
wire w0;    //: /sn:0 /dp:1 {0}(1071,316)(1058,316)(1058,280)(1044,280){1}
wire w20;    //: /sn:0 {0}(1096,396)(1112,396)(1112,366)(1150,366){1}
wire w30;    //: /sn:0 {0}(380,233)(380,184){1}
//: {2}(382,182)(446,182){3}
//: {4}(450,182)(507,182){5}
//: {6}(511,182)(663,182){7}
//: {8}(509,184)(509,231){9}
//: {10}(448,184)(448,231){11}
//: {12}(378,182)(312,182){13}
//: {14}(310,180)(310,124){15}
//: {16}(308,182)(242,182){17}
//: {18}(238,182)(191,182){19}
//: {20}(240,184)(240,231){21}
//: {22}(310,184)(310,233){23}
wire w18;    //: /sn:0 {0}(1047,410)(1059,410)(1059,398)(1075,398){1}
wire w19;    //: /sn:0 {0}(871,379)(871,391)(878,391){1}
//: {2}(880,389)(880,355){3}
//: {4}(882,353)(1071,353){5}
//: {6}(880,351)(880,321){7}
//: {8}(882,319)(1023,319){9}
//: {10}(880,317)(880,280)(1023,280){11}
//: {12}(880,393)(880,463){13}
wire w10;    //: /sn:0 {0}(1023,275)(860,275)(860,312){1}
//: {2}(862,314)(1023,314){3}
//: {4}(860,316)(860,387){5}
//: {6}(858,389)(850,389)(850,379){7}
//: {8}(860,391)(860,405){9}
//: {10}(862,407)(1026,407){11}
//: {12}(860,409)(860,463){13}
wire w1;    //: /sn:0 {0}(1023,324)(898,324)(898,463){1}
wire w32;    //: /sn:0 {0}(370,233)(370,164){1}
//: {2}(372,162)(436,162){3}
//: {4}(440,162)(497,162){5}
//: {6}(501,162)(665,162){7}
//: {8}(499,164)(499,231){9}
//: {10}(438,164)(438,231){11}
//: {12}(368,162)(302,162){13}
//: {14}(300,160)(300,124){15}
//: {16}(298,162)(232,162){17}
//: {18}(228,162)(191,162){19}
//: {20}(230,164)(230,231){21}
//: {22}(300,164)(300,233){23}
wire w41;    //: /sn:0 {0}(494,231)(494,154){1}
//: {2}(496,152)(665,152){3}
//: {4}(492,152)(435,152){5}
//: {6}(431,152)(367,152){7}
//: {8}(363,152)(297,152){9}
//: {10}(295,150)(295,124){11}
//: {12}(293,152)(227,152){13}
//: {14}(223,152)(191,152){15}
//: {16}(225,154)(225,231){17}
//: {18}(295,154)(295,233){19}
//: {20}(365,154)(365,233){21}
//: {22}(433,154)(433,231){23}
wire w15;    //: /sn:0 {0}(1044,321)(1071,321){1}
wire w5;    //: /sn:0 {0}(191,192)(243,192){1}
//: {2}(247,192)(313,192){3}
//: {4}(317,192)(383,192){5}
//: {6}(387,192)(451,192){7}
//: {8}(455,192)(512,192){9}
//: {10}(516,192)(665,192){11}
//: {12}(514,194)(514,231){13}
//: {14}(453,194)(453,231){15}
//: {16}(385,194)(385,233){17}
//: {18}(315,190)(315,124){19}
//: {20}(315,194)(315,233){21}
//: {22}(245,194)(245,231){23}
wire w9;    //: /sn:0 /dp:1 {0}(1023,270)(840,270)(840,307){1}
//: {2}(842,309)(1023,309){3}
//: {4}(840,311)(840,386){5}
//: {6}(838,388)(825,388)(825,381){7}
//: {8}(840,390)(840,463){9}
//: enddecls

  and g4 (.I0(w7), .I1(!w5), .I2(w30), .I3(!w39), .I4(w32), .I5(w41), .Z(MemWrite));   //: @(378,244) /sn:0 /R:3 /w:[ 17 17 0 21 0 21 5 ]
  //: comment g8 /dolink:0 /link:"" @(275,235) /sn:0 /R:3
  //: /line:"lw"
  //: /end
  //: output g44 (Jump) @(568,320) /sn:0 /w:[ 0 ]
  //: joint g75 (w10) @(860, 407) /w:[ 10 9 -1 12 ]
  and g3 (.I0(w7), .I1(!w5), .I2(!w30), .I3(!w39), .I4(w32), .I5(w41), .Z(MemToReg));   //: @(308,244) /sn:0 /R:3 /w:[ 21 21 23 19 23 19 5 ]
  //: joint g16 (w41) @(494, 152) /w:[ 2 -1 4 1 ]
  //: output g47 (MemWrite) @(568,423) /sn:0 /w:[ 0 ]
  //: joint g17 (w39) @(235, 172) /w:[ 13 -1 14 16 ]
  //: joint g26 (w30) @(448, 182) /w:[ 4 -1 3 10 ]
  led g90 (.I(Branch));   //: @(923,458) /sn:0 /w:[ 11 ] /type:0
  led g109 (.I(funct));   //: @(811,417) /sn:0 /R:1 /w:[ 11 ] /type:2
  and g2 (.I0(!w7), .I1(!w5), .I2(!w30), .I3(!w39), .I4(!w32), .I5(!w41), .Z(RegDst));   //: @(238,242) /sn:0 /R:3 /w:[ 0 23 21 17 21 17 25 ]
  //: joint g23 (w7) @(519, 202) /w:[ 10 -1 9 12 ]
  //: joint g30 (w32) @(230, 162) /w:[ 17 -1 18 20 ]
  //: joint g74 (RegDst) @(957, 412) /w:[ 10 9 -1 12 ]
  //: joint g91 (Branch) @(934, 478) /w:[ -1 9 10 12 ]
  led g92 (.I(RegDst));   //: @(215,263) /sn:0 /w:[ 27 ] /type:0
  tran g86(.Z(w1), .I(funct[3]));   //: @(898,466) /sn:0 /R:1 /w:[ 1 2 1 ] /ss:0
  concat g1 (.I0(w41), .I1(w32), .I2(w39), .I3(w30), .I4(w5), .I5(w7), .Z(op));   //: @(186,177) /sn:0 /R:2 /w:[ 15 19 15 19 0 23 1 ] /dr:0
  //: joint g24 (w30) @(509, 182) /w:[ 6 -1 5 8 ]
  //: joint g39 (w30) @(380, 182) /w:[ 2 -1 12 1 ]
  //: joint g77 (Branch) @(934, 393) /w:[ 1 2 -1 8 ]
  //: joint g104 (w9) @(840, 388) /w:[ -1 5 6 8 ]
  //: comment g111 /dolink:0 /link:"" @(1025,418) /sn:0
  //: /line:"sub/slt"
  //: /end
  //: joint g29 (w32) @(438, 162) /w:[ 4 -1 3 10 ]
  //: frame g60 @(92,47) /sn:0 /wi:629 /ht:506 /tx:"Unitat Control"
  //: joint g110 (funct) @(824, 468) /w:[ 9 10 12 -1 ]
  or g51 (.I0(MemWrite), .I1(MemToReg), .Z(ALUSrc));   //: @(536,444) /sn:0 /w:[ 9 11 1 ]
  //: joint g18 (w39) @(305, 172) /w:[ 9 10 12 18 ]
  //: comment g70 /dolink:0 /link:"" @(904,429) /sn:0 /R:2
  //: /line:"op0"
  //: /end
  //: joint g82 (w9) @(840, 309) /w:[ 2 1 -1 4 ]
  //: comment g10 /dolink:0 /link:"" @(409,239) /sn:0 /R:3
  //: /line:"beq"
  //: /end
  //: joint g25 (w32) @(499, 162) /w:[ 6 -1 5 8 ]
  tran g65(.Z(w9), .I(funct[0]));   //: @(840,466) /sn:0 /R:1 /w:[ 9 8 7 ] /ss:0
  //: joint g94 (MemToReg) @(308, 285) /w:[ -1 4 6 3 ]
  led g103 (.I(w9));   //: @(825,374) /sn:0 /w:[ 7 ] /type:0
  //: output g64 (ALUOp) @(1188,361) /sn:0 /w:[ 3 ]
  led g107 (.I(w19));   //: @(871,372) /sn:0 /w:[ 0 ] /type:0
  //: joint g72 (RegDst) @(957, 358) /w:[ 6 5 -1 8 ]
  //: output g49 (ALUSrc) @(568,444) /sn:0 /w:[ 0 ]
  and g6 (.I0(!w7), .I1(!w5), .I2(!w30), .I3(!w39), .I4(w32), .I5(!w41), .Z(Jump));   //: @(507,242) /sn:0 /R:3 /w:[ 13 13 9 0 9 0 3 ]
  //: output g50 (RegWrite) @(569,468) /sn:0 /w:[ 1 ]
  //: comment g7 /dolink:0 /link:"" @(175,236) /sn:0 /R:3
  //: /line:"Tipus R"
  //: /end
  //: comment g9 /dolink:0 /link:"" @(345,235) /sn:0 /R:3
  //: /line:"sw"
  //: /end
  //: joint g35 (w5) @(315, 192) /w:[ 4 18 3 20 ]
  //: output g56 (MemRead) @(567,371) /sn:0 /w:[ 1 ]
  //: joint g58 (MemWrite) @(378, 423) /w:[ 1 2 -1 8 ]
  tran g68(.Z(w10), .I(funct[1]));   //: @(860,466) /sn:0 /R:1 /w:[ 13 6 5 ] /ss:0
  or g73 (.I0(Branch), .I1(w18), .Z(w20));   //: @(1086,396) /sn:0 /w:[ 0 1 0 ]
  //: joint g22 (w5) @(514, 192) /w:[ 10 -1 9 12 ]
  //: joint g31 (w30) @(240, 182) /w:[ 17 -1 18 20 ]
  //: joint g59 (MemToReg) @(308, 446) /w:[ 10 9 -1 12 ]
  or g71 (.I0(w0), .I1(w15), .Z(w6));   //: @(1082,319) /sn:0 /w:[ 0 1 0 ]
  //: joint g98 (Branch) @(446, 281) /w:[ -1 18 20 17 ]
  //: joint g102 (ALUOp) @(1170, 361) /w:[ 2 -1 1 4 ]
  //: joint g85 (RegDst) @(957, 334) /w:[ 1 2 -1 4 ]
  concat g67 (.I0(w6), .I1(w4), .I2(w20), .I3(w3), .Z(ALUOp));   //: @(1155,361) /sn:0 /w:[ 1 1 1 0 0 ] /dr:1
  //: frame g87 @(753,244) /sn:0 /wi:510 /ht:308 /tx:"ALU Control"
  //: joint g83 (w10) @(860, 314) /w:[ 2 1 -1 4 ]
  led g99 (.I(Jump));   //: @(486,267) /sn:0 /w:[ 5 ] /type:0
  //: joint g33 (w7) @(250, 202) /w:[ 2 -1 22 1 ]
  //: joint g36 (w30) @(310, 182) /w:[ 13 14 16 22 ]
  //: joint g41 (w5) @(385, 192) /w:[ 6 -1 5 16 ]
  //: output g45 (Branch) @(567,345) /sn:0 /w:[ 15 ]
  and g54 (.I0(w41), .I1(w32), .I2(!w39), .I3(!w30), .I4(!w5), .I5(w7), .Z(MemRead));   //: @(307,113) /sn:0 /R:1 /w:[ 11 15 11 15 19 19 0 ]
  //: joint g40 (w7) @(390, 202) /w:[ 6 -1 5 16 ]
  //: comment g42 /dolink:0 /link:"" @(791,48) /sn:0 /R:3
  //: /line:"         opcode      func      ALUOp   ALUCtrl"
  //: /line:"add     00 0000     10 0000     10      0010"
  //: /line:"sub     00 0000     10 0010     10      0110"
  //: /line:"and     00 0000     10 0100     10      0000"
  //: /line:"or      00 0000     10 0101     10      0001"
  //: /line:"slt     00 0000     10 1010     10      0111"
  //: /line:""
  //: /line:"lw      10 0011     XX XXXX     00      0010"
  //: /line:"sw      10 1011     XX XXXX     00      0010"
  //: /line:"beq     00 0100     XX XXXX     01      0110"
  //: /line:"j       00 0010     XX XXXX     XX      XXXX"
  //: /end
  or g52 (.I0(MemToReg), .I1(RegDst), .Z(RegWrite));   //: @(535,468) /sn:0 /w:[ 13 19 0 ]
  tran g69(.Z(w19), .I(funct[2]));   //: @(880,466) /sn:0 /R:1 /w:[ 13 4 3 ] /ss:0
  and g81 (.I0(!w9), .I1(w10), .I2(!w19), .I3(w1), .I4(!Branch), .I5(RegDst), .Z(w15));   //: @(1034,321) /sn:0 /w:[ 3 3 9 0 5 0 0 ]
  //: supply0 g66 (w3) @(1129,399) /sn:0 /w:[ 1 ]
  //: joint g12 (w41) @(225, 152) /w:[ 13 -1 14 16 ]
  //: joint g108 (w19) @(880, 391) /w:[ -1 2 1 12 ]
  //: joint g28 (w7) @(458, 202) /w:[ 8 -1 7 14 ]
  //: joint g34 (w7) @(320, 202) /w:[ 4 18 3 20 ]
  //: output g46 (MemToReg) @(567,392) /sn:0 /w:[ 0 ]
  //: comment g57 /dolink:0 /link:"" @(357,73) /sn:0
  //: /line:"1 cable no pot conectarse a 2 sortides"
  //: /line:"Buffer A=4u R=4T"
  //: /line:"AND2 A=6u R=6T"
  //: /line:"Sacrificar 2 de area per 0 Retard (en paralel)"
  //: /end
  //: joint g106 (w10) @(860, 389) /w:[ -1 5 6 8 ]
  and g5 (.I0(!w7), .I1(!w5), .I2(!w30), .I3(w39), .I4(!w32), .I5(!w41), .Z(Branch));   //: @(446,242) /sn:0 /R:3 /w:[ 15 15 11 23 11 23 19 ]
  //: comment g11 /dolink:0 /link:"" @(480,241) /sn:0 /R:3
  //: /line:"j"
  //: /end
  //: joint g14 (w41) @(365, 152) /w:[ 7 -1 8 20 ]
  //: joint g84 (w19) @(880, 319) /w:[ 8 10 -1 7 ]
  //: comment g112 /dolink:0 /link:"" @(1083,402) /sn:0
  //: /line:"beq"
  //: /end
  //: joint g96 (MemWrite) @(378, 283) /w:[ -1 4 6 3 ]
  nand g114 (.I0(w19), .I1(RegDst), .Z(w4));   //: @(1082,356) /sn:0 /w:[ 5 7 0 ]
  //: joint g19 (w39) @(375, 172) /w:[ 7 -1 8 20 ]
  //: joint g21 (w39) @(504, 172) /w:[ 2 -1 4 1 ]
  //: joint g61 (Branch) @(446, 345) /w:[ 14 16 -1 13 ]
  //: joint g79 (Branch) @(934, 329) /w:[ 4 6 -1 3 ]
  //: joint g78 (w19) @(880, 353) /w:[ 4 6 -1 3 ]
  //: joint g20 (w39) @(443, 172) /w:[ 5 -1 6 22 ]
  //: joint g32 (w5) @(245, 192) /w:[ 2 -1 1 22 ]
  //: comment g113 /dolink:0 /link:"" @(1018,362) /sn:0
  //: /line:"NOT and/or"
  //: /end
  //: input g63 (funct) @(807,468) /sn:0 /w:[ 13 ]
  led g93 (.I(MemToReg));   //: @(294,267) /sn:0 /w:[ 7 ] /type:0
  led g97 (.I(Branch));   //: @(417,266) /sn:0 /w:[ 21 ] /type:0
  //: joint g100 (Jump) @(507, 282) /w:[ -1 2 4 1 ]
  led g105 (.I(w10));   //: @(850,372) /sn:0 /w:[ 7 ] /type:0
  //: input g0 (op) @(147,177) /sn:0 /w:[ 0 ]
  //: joint g15 (w41) @(433, 152) /w:[ 5 -1 6 22 ]
  //: joint g38 (w32) @(370, 162) /w:[ 2 -1 12 1 ]
  //: output g43 (RegDst) @(567,294) /sn:0 /w:[ 23 ]
  //: joint g89 (RegDst) @(957, 479) /w:[ 14 13 -1 16 ]
  led g101 (.I(ALUOp));   //: @(1170,399) /sn:0 /R:2 /w:[ 5 ] /type:2
  //: joint g27 (w5) @(453, 192) /w:[ 8 -1 7 14 ]
  //: joint g48 (MemToReg) @(308, 392) /w:[ 1 2 -1 8 ]
  //: joint g37 (w32) @(300, 162) /w:[ 13 14 16 22 ]
  //: comment g62 /dolink:0 /link:"" @(964,428) /sn:0 /R:2
  //: /line:"op1"
  //: /end
  //: joint g55 (RegDst) @(238, 470) /w:[ 18 20 -1 17 ]
  and g80 (.I0(w9), .I1(!w10), .I2(w19), .I3(!Branch), .I4(RegDst), .Z(w0));   //: @(1034,280) /sn:0 /w:[ 0 0 11 7 3 1 ]
  led g88 (.I(RegDst));   //: @(974,464) /sn:0 /w:[ 15 ] /type:0
  led g95 (.I(MemWrite));   //: @(362,268) /sn:0 /w:[ 7 ] /type:0
  //: joint g13 (w41) @(295, 152) /w:[ 9 10 12 18 ]
  //: joint g53 (RegDst) @(238, 294) /w:[ 22 24 26 21 ]
  and g76 (.I0(w10), .I1(RegDst), .Z(w18));   //: @(1037,410) /sn:0 /w:[ 11 11 0 ]

endmodule

module main;    //: root_module
wire [5:0] w4;    //: /sn:0 /dp:1 {0}(668,48)(693,48){1}
wire w3;    //: /sn:0 {0}(843,19)(892,19){1}
wire w29;    //: /sn:0 {0}(843,-73)(893,-73){1}
wire w30;    //: /sn:0 {0}(843,-96)(893,-96){1}
wire w23;    //: /sn:0 /dp:1 {0}(843,-50)(893,-50){1}
wire [3:0] SignExtOut;    //: /sn:0 /dp:1 {0}(933,-2)(921,-2){1}
//: {2}(917,-2)(843,-2){3}
//: {4}(919,0)(919,35)(1031,35)(1031,20){5}
wire w31;    //: /sn:0 {0}(843,-116)(892,-116){1}
wire w8;    //: /sn:0 /dp:1 {0}(843,62)(892,62){1}
wire w27;    //: /sn:0 {0}(843,-24)(893,-24){1}
wire [5:0] w5;    //: /sn:0 /dp:1 {0}(668,3)(693,3){1}
wire w9;    //: /sn:0 {0}(843,35)(893,35){1}
//: enddecls

  //: joint g3 (SignExtOut) @(919, -2) /w:[ 1 -1 2 4 ]
  led g26 (.I(w29));   //: @(900,-73) /sn:0 /R:3 /w:[ 1 ] /type:0
  led g2 (.I(SignExtOut));   //: @(1031,13) /sn:0 /w:[ 5 ] /type:1
  led g23 (.I(w30));   //: @(900,-96) /sn:0 /R:3 /w:[ 1 ] /type:0
  led g30 (.I(w27));   //: @(900,-24) /sn:0 /R:3 /w:[ 1 ] /type:0
  //: dip g1 (w5) @(630,3) /sn:0 /R:1 /w:[ 0 ] /st:2
  led g29 (.I(w23));   //: @(900,-50) /sn:0 /R:3 /w:[ 1 ] /type:0
  led g31 (.I(w3));   //: @(899,19) /sn:0 /R:3 /w:[ 1 ] /type:0
  led g33 (.I(w9));   //: @(900,35) /sn:0 /R:3 /w:[ 1 ] /type:0
  led g81 (.I(SignExtOut));   //: @(940,-2) /sn:0 /R:3 /w:[ 0 ] /type:2
  led g21 (.I(w31));   //: @(899,-116) /sn:0 /R:3 /w:[ 1 ] /type:0
  //: dip g0 (w4) @(630,48) /sn:0 /R:1 /w:[ 0 ] /st:33
  CONTROL g38 (.funct(w4), .op(w5), .MemWrite(w3), .RegDst(w31), .Jump(w30), .Branch(w29), .MemRead(w23), .MemToReg(w27), .ALUOp(SignExtOut), .ALUSrc(w9), .RegWrite(w8));   //: @(694, -139) /sz:(148, 230) /sn:0 /p:[ Li0>1 Li1>1 Ro0<0 Ro1<0 Ro2<0 Ro3<0 Ro4<0 Ro5<0 Ro6<3 Ro7<0 Ro8<0 ]
  led g37 (.I(w8));   //: @(899,62) /sn:0 /R:3 /w:[ 1 ] /type:0

endmodule
