//: version "1.8.7"

module Zero(o, i);
//: interface  /sz:(40, 40) /bd:[ Li0>i[31:0](21/40) Ro0<o(22/40) ]
input [31:0] i;    //: /sn:0 {0}(441,304)(494,304){1}
output o;    //: /sn:0 /dp:1 {0}(645,292)(645,317)(802,317){1}
wire w0;    //: /sn:0 {0}(632,194)(645,194)(645,244){1}
wire [31:0] w1;    //: /sn:0 /dp:1 {0}(496,228)(496,252)(631,252){1}
wire [31:0] w5;    //: /sn:0 /dp:1 {0}(660,268)(787,268)(787,239){1}
wire [31:0] w9;    //: /sn:0 {0}(568,303)(602,303)(602,284)(631,284){1}
//: enddecls

  led g4 (.I(w5));   //: @(787,232) /sn:0 /w:[ 1 ] /type:3
  //: dip g3 (w1) @(496,218) /sn:0 /w:[ 0 ] /st:0
  //: switch g2 (w0) @(615,194) /sn:0 /w:[ 0 ] /st:0
  //: output g1 (o) @(799,317) /sn:0 /w:[ 1 ]
  Ca2 g6 (.in(i), .out(w9));   //: @(495, 282) /sz:(72, 40) /sn:0 /p:[ Li0>1 Ro0<0 ]
  add g5 (.A(w9), .B(w1), .S(w5), .CI(w0), .CO(o));   //: @(647,268) /sn:0 /R:1 /w:[ 1 1 0 1 0 ]
  //: input g0 (i) @(439,304) /sn:0 /w:[ 0 ]

endmodule

module SignExtend(D32b, D16b);
//: interface  /sz:(207, 73) /bd:[ Li0>D16b[15:0](37/73) Ro0<D32b[31:0](36/73) ]
output [31:0] D32b;    //: /sn:0 /dp:1 {0}(737,171)(678,171)(678,167)(641,167){1}
supply0 [15:0] w0;    //: /sn:0 {0}(153,107)(153,98)(169,98)(169,162)(635,162){1}
input [15:0] D16b;    //: /sn:0 /dp:1 {0}(635,172)(149,172){1}
//: enddecls

  //: output g3 (D32b) @(734,171) /sn:0 /w:[ 0 ]
  concat g2 (.I0(D16b), .I1(w0), .Z(D32b));   //: @(640,167) /sn:0 /w:[ 0 1 1 ] /dr:0
  //: supply0 g1 (w0) @(153,113) /sn:0 /w:[ 0 ]
  //: input g0 (D16b) @(147,172) /sn:0 /w:[ 1 ]

endmodule

module Ca2(out, in);
//: interface  /sz:(72, 40) /bd:[ Li0>in[31:0](22/40) Ro0<out[31:0](21/40) ]
input [31:0] in;    //: /sn:0 {0}(494,347)(552,347){1}
supply0 w0;    //: /sn:0 {0}(551,307)(551,297)(566,297)(566,339){1}
output [31:0] out;    //: /sn:0 /dp:1 {0}(581,363)(639,363){1}
wire [31:0] w1;    //: /sn:0 /dp:1 {0}(484,393)(484,379)(552,379){1}
wire w2;    //: /sn:0 /dp:1 {0}(581,419)(581,429)(566,429)(566,387){1}
//: enddecls

  //: supply0 g4 (w0) @(551,313) /sn:0 /w:[ 0 ]
  //: dip g3 (w1) @(484,404) /sn:0 /R:2 /w:[ 0 ] /st:1
  add g2 (.A(w1), .B(in), .S(out), .CI(w0), .CO(w2));   //: @(568,363) /sn:0 /R:1 /w:[ 1 1 0 1 1 ]
  //: output g1 (out) @(636,363) /sn:0 /w:[ 1 ]
  led g5 (.I(w2));   //: @(581,412) /sn:0 /w:[ 0 ] /type:0
  //: input g0 (in) @(492,347) /sn:0 /w:[ 0 ]

endmodule

module ALU(Result, Zero, B, A, ALU_OP);
//: interface  /sz:(94, 87) /bd:[ Ti0>ALU_OP[3:0](45/94) Li0>B[31:0](70/87) Li1>A[31:0](30/87) Ro0<Result[31:0](66/87) Ro1<Zero(32/87) ]
input [31:0] B;    //: /sn:0 /dp:1 {0}(571,193)(270,193)(270,280){1}
//: {2}(272,282)(576,282){3}
//: {4}(270,284)(270,358){5}
//: {6}(268,360)(131,360)(131,153){7}
//: {8}(270,362)(270,411){9}
//: {10}(268,413)(222,413){11}
//: {12}(270,415)(270,454){13}
//: {14}(272,456)(569,456){15}
//: {16}(270,458)(270,599)(446,599){17}
output Zero;    //: /sn:0 {0}(1411,566)(1505,566){1}
input [31:0] A;    //: /sn:0 {0}(317,322)(359,322){1}
//: {2}(361,320)(361,279){3}
//: {4}(363,277)(576,277){5}
//: {6}(361,275)(361,188)(571,188){7}
//: {8}(361,324)(361,344){9}
//: {10}(363,346)(513,346)(513,112){11}
//: {12}(361,348)(361,422){13}
//: {14}(363,424)(569,424){15}
//: {16}(361,426)(361,566)(570,566){17}
output [31:0] Result;    //: /sn:0 /dp:1 {0}(1084,348)(1317,348){1}
//: {2}(1321,348)(1415,348){3}
//: {4}(1319,350)(1319,565)(1369,565){5}
input [3:0] ALU_OP;    //: /sn:0 /dp:1 {0}(1071,325)(1071,123)(1007,123){1}
wire [31:0] w6;    //: /sn:0 /dp:1 {0}(1021,699)(1021,561){1}
wire [31:0] w13;    //: /sn:0 {0}(1011,532)(1011,503){1}
//: {2}(1013,501)(1162,501)(1162,493){3}
//: {4}(1011,499)(1011,346)(1055,346){5}
wire w16;    //: /sn:0 {0}(584,606)(584,636)(610,636)(610,626){1}
wire [31:0] w3;    //: /sn:0 /dp:1 {0}(1055,328)(710,328)(710,440)(658,440){1}
//: {2}(654,440)(598,440){3}
//: {4}(656,442)(656,476)(801,476)(801,536)(855,536)(855,704)(681,704)(681,694){5}
wire w22;    //: /sn:0 {0}(545,525)(584,525)(584,558){1}
wire [31:0] w0;    //: /sn:0 {0}(520,598)(570,598){1}
wire [31:0] w20;    //: /sn:0 {0}(953,644)(953,607)(964,607){1}
//: {2}(968,607)(1001,607)(1001,561){3}
//: {4}(966,605)(966,468)(956,468){5}
//: {6}(954,466)(954,374)(1055,374){7}
//: {8}(952,468)(940,468){9}
//: {10}(938,466)(938,370)(1055,370){11}
//: {12}(936,468)(922,468){13}
//: {14}(920,466)(920,367)(1055,367){15}
//: {16}(918,468)(903,468){17}
//: {18}(901,466)(901,363)(1055,363){19}
//: {20}(899,468)(882,468){21}
//: {22}(880,466)(880,360)(1055,360){23}
//: {24}(878,468)(864,468){25}
//: {26}(862,466)(862,356)(1055,356){27}
//: {28}(860,468)(838,468){29}
//: {30}(836,466)(836,353)(1055,353){31}
//: {32}(834,468)(813,468){33}
//: {34}(811,466)(811,349)(1055,349){35}
//: {36}(809,468)(794,468){37}
//: {38}(792,466)(792,339)(1055,339){39}
//: {40}(790,468)(770,468){41}
//: {42}(768,466)(768,335)(1055,335){43}
//: {44}(766,468)(732,468)(732,332)(1055,332){45}
wire w23;    //: /sn:0 {0}(537,372)(583,372)(583,416){1}
wire w21;    //: /sn:0 {0}(583,464)(583,498)(600,498)(600,488){1}
wire [31:0] w1;    //: /sn:0 /dp:1 {0}(1055,321)(716,321)(716,191)(592,191){1}
wire w11;    //: /sn:0 {0}(697,545)(988,545){1}
wire [31:0] w2;    //: /sn:0 /dp:1 {0}(1055,325)(689,325)(689,280)(597,280){1}
wire [31:0] w9;    //: /sn:0 /dp:3 {0}(599,582)(693,582)(693,545){1}
//: {2}(693,544)(693,342)(1055,342){3}
//: enddecls

  add g8 (.A(w0), .B(A), .S(w9), .CI(w22), .CO(w16));   //: @(586,582) /sn:0 /R:1 /w:[ 1 17 0 1 0 ]
  //: output g4 (Result) @(1412,348) /sn:0 /w:[ 3 ]
  led g44 (.I(A));   //: @(513,105) /sn:0 /w:[ 11 ] /type:3
  //: joint g16 (B) @(270, 282) /w:[ 2 1 -1 4 ]
  //: output g3 (Zero) @(1502,566) /sn:0 /w:[ 1 ]
  //: joint g47 (w3) @(656, 440) /w:[ 1 -1 2 4 ]
  led g26 (.I(w13));   //: @(1162,486) /sn:0 /w:[ 3 ] /type:3
  //: joint g17 (B) @(270, 413) /w:[ -1 9 10 12 ]
  //: input g2 (B) @(220,413) /sn:0 /w:[ 11 ]
  //: joint g30 (Result) @(1319, 348) /w:[ 2 -1 1 4 ]
  //: comment g23 /dolink:0 /link:"" @(1052,527) /sn:0
  //: /line:"if (A < B)   // bit 31 = 1"
  //: /line:"   ALU = 1;"
  //: /line:"else         // bit 31 = 0"
  //: /line:"   ALU = 0;"
  //: /end
  //: joint g39 (w20) @(811, 468) /w:[ 33 34 36 -1 ]
  //: dip g24 (w6) @(1021,710) /sn:0 /R:2 /w:[ 0 ] /st:1
  //: input g1 (A) @(315,322) /sn:0 /w:[ 0 ]
  Zero g29 (.i(Result), .o(Zero));   //: @(1370, 544) /sz:(40, 40) /sn:0 /p:[ Li0>5 Ro0<0 ]
  //: joint g18 (B) @(270, 456) /w:[ 14 13 -1 16 ]
  //: dip g25 (w20) @(953,655) /sn:0 /R:2 /w:[ 0 ] /st:0
  //: switch g10 (w22) @(528,525) /sn:0 /w:[ 0 ] /st:0
  or g6 (.I0(A), .I1(B), .Z(w2));   //: @(587,280) /sn:0 /w:[ 5 3 1 ]
  //: joint g35 (w20) @(901, 468) /w:[ 17 18 20 -1 ]
  mux g7 (.I0(w1), .I1(w2), .I2(w3), .I3(w20), .I4(w20), .I5(w20), .I6(w9), .I7(w13), .I8(w20), .I9(w20), .I10(w20), .I11(w20), .I12(w20), .I13(w20), .I14(w20), .I15(w20), .S(ALU_OP), .Z(Result));   //: @(1071,348) /sn:0 /R:1 /w:[ 0 0 0 45 43 39 3 5 35 31 27 23 19 15 11 7 0 0 ] /ss:1 /do:1
  add g9 (.A(B), .B(A), .S(w3), .CI(w23), .CO(w21));   //: @(585,440) /sn:0 /R:1 /w:[ 15 15 3 1 0 ]
  //: joint g31 (w20) @(966, 607) /w:[ 2 4 1 -1 ]
  tran g22(.Z(w11), .I(w9[31]));   //: @(691,545) /sn:0 /R:2 /w:[ 0 1 2 ] /ss:1
  //: joint g41 (w20) @(768, 468) /w:[ 41 42 44 -1 ]
  //: joint g36 (w20) @(880, 468) /w:[ 21 22 24 -1 ]
  //: joint g33 (w20) @(938, 468) /w:[ 9 10 12 -1 ]
  //: joint g45 (A) @(361, 346) /w:[ 10 9 -1 12 ]
  //: joint g40 (w20) @(792, 468) /w:[ 37 38 40 -1 ]
  led g42 (.I(B));   //: @(131,146) /sn:0 /w:[ 7 ] /type:3
  //: input g12 (ALU_OP) @(1005,123) /sn:0 /w:[ 1 ]
  //: joint g34 (w20) @(920, 468) /w:[ 13 14 16 -1 ]
  //: comment g28 /dolink:0 /link:"" @(845,478) /sn:0
  //: /line:"not used pins"
  //: /line:""
  //: /end
  led g46 (.I(w3));   //: @(681,687) /sn:0 /w:[ 5 ] /type:3
  //: joint g14 (A) @(361, 322) /w:[ -1 2 1 8 ]
  //: switch g11 (w23) @(520,372) /sn:0 /w:[ 0 ] /st:0
  and g5 (.I0(A), .I1(B), .Z(w1));   //: @(582,191) /sn:0 /w:[ 7 0 1 ]
  mux g21 (.I0(w20), .I1(w6), .S(w11), .Z(w13));   //: @(1011,545) /sn:0 /R:2 /w:[ 3 1 1 0 ] /ss:1 /do:1
  led g19 (.I(w16));   //: @(610,619) /sn:0 /w:[ 1 ] /type:0
  led g20 (.I(w21));   //: @(600,481) /sn:0 /w:[ 1 ] /type:0
  //: joint g32 (w20) @(954, 468) /w:[ 5 6 8 -1 ]
  //: joint g38 (w20) @(836, 468) /w:[ 29 30 32 -1 ]
  //: joint g15 (A) @(361, 424) /w:[ 14 13 -1 16 ]
  Ca2 g0 (.in(B), .out(w0));   //: @(447, 577) /sz:(72, 40) /sn:0 /p:[ Li0>17 Ro0<0 ]
  //: joint g43 (B) @(270, 360) /w:[ -1 5 6 8 ]
  //: joint g27 (w13) @(1011, 501) /w:[ 2 4 -1 1 ]
  //: joint g37 (w20) @(862, 468) /w:[ 25 26 28 -1 ]
  //: joint g13 (A) @(361, 277) /w:[ 4 6 -1 3 ]

endmodule

module BRegs32x32(Read2, Write, Read1, Data2, Data1, clr, clk, RegWrite, WriteData);
//: interface  /sz:(147, 182) /bd:[ Ti0>clr(66/147) Li0>Read1[4:0](32/182) Li1>Read2[4:0](72/182) Li2>Write[4:0](108/182) Li3>WriteData[31:0](148/182) Bi0>clk(108/147) Bi1>RegWrite(40/147) Ro0<Data1[31:0](47/182) Ro1<Data2[31:0](139/182) ]
output [31:0] Data2;    //: /sn:0 {0}(668,485)(668,472)(669,472)(669,445){1}
input [4:0] Write;    //: /sn:0 {0}(-238,-38)(-138,-38)(-138,-37)(-66,-37){1}
//: {2}(-65,-37)(-28,-37){3}
//: {4}(-27,-37)(-16,-37){5}
input [31:0] WriteData;    //: /sn:0 {0}(669,157)(669,75)(481,75){1}
//: {2}(477,75)(292,75){3}
//: {4}(288,75)(89,75){5}
//: {6}(85,75)(-104,75)(-104,73)(-237,73){7}
//: {8}(87,77)(87,157){9}
//: {10}(290,77)(290,107)(291,107)(291,152){11}
//: {12}(479,77)(479,157){13}
output [31:0] Data1;    //: /sn:0 {0}(59,382)(59,465){1}
supply1 w21;    //: /sn:0 {0}(82,3)(57,3)(57,-11){1}
input clr;    //: /sn:0 {0}(721,193)(731,193)(731,-83)(543,-83){1}
//: {2}(539,-83)(355,-83){3}
//: {4}(351,-83)(150,-83){5}
//: {6}(146,-83)(-44,-83)(-44,-92)(-235,-92){7}
//: {8}(148,-81)(148,193)(139,193){9}
//: {10}(353,-81)(353,188)(343,188){11}
//: {12}(541,-81)(541,193)(531,193){13}
input RegWrite;    //: /sn:0 {0}(-237,263)(-71,263){1}
//: {2}(-67,263)(171,263){3}
//: {4}(175,263)(370,263){5}
//: {6}(374,263)(552,263)(552,219)(556,219){7}
//: {8}(372,261)(372,219)(383,219){9}
//: {10}(173,261)(173,214)(183,214){11}
//: {12}(-69,261)(-69,219)(-38,219){13}
input clk;    //: /sn:0 {0}(556,214)(542,214)(542,285)(364,285){1}
//: {2}(362,283)(362,214)(383,214){3}
//: {4}(360,285)(167,285){5}
//: {6}(165,283)(165,209)(183,209){7}
//: {8}(163,285)(-56,285){9}
//: {10}(-58,283)(-58,214)(-38,214){11}
//: {12}(-60,285)(-237,285){13}
input [4:0] Read1;    //: {0}(-237,96)(-208,96)(-208,95)(-124,95){1}
//: {2}(-123,95)(-96,95){3}
//: {4}(-95,95)(-78,95){5}
input [4:0] Read2;    //: {0}(-237,145)(-141,145){1}
//: {2}(-140,145)(-123,145)(-123,144)(-94,144){3}
//: {4}(-93,144)(-79,144){5}
wire [1:0] w6;    //: /sn:0 {0}(36,369)(-123,369)(-123,99){1}
wire w16;    //: /sn:0 {0}(39,205)(-50,205)(-50,39)(88,39)(88,19){1}
wire w4;    //: /sn:0 {0}(112,19)(112,46)(370,46)(370,205)(431,205){1}
wire [31:0] w3;    //: /sn:0 {0}(77,353)(77,334)(659,334)(659,228){1}
wire [31:0] R2;    //: {0}(65,353)(65,319)(469,319)(469,228){1}
wire [31:0] w0;    //: /sn:0 {0}(651,416)(651,398)(105,398)(105,228){1}
wire w22;    //: /sn:0 {0}(404,217)(431,217){1}
wire w20;    //: /sn:0 {0}(124,19)(124,29)(556,29)(556,205)(621,205){1}
wire [2:0] w19;    //: /sn:0 {0}(431,169)(419,169)(419,109){1}
//: {2}(421,107)(606,107)(606,169)(621,169){3}
//: {4}(417,107)(297,107)(297,106)(231,106){5}
//: {6}(227,106)(25,106){7}
//: {8}(21,106)(-95,106)(-95,99){9}
//: {10}(23,108)(23,169)(39,169){11}
//: {12}(229,108)(229,164)(243,164){13}
wire [2:0] w18;    //: /sn:0 {0}(431,180)(402,180)(402,125){1}
//: {2}(404,123)(589,123)(589,180)(621,180){3}
//: {4}(400,123)(279,123)(279,122)(212,122){5}
//: {6}(208,122)(8,122){7}
//: {8}(4,122)(-93,122)(-93,139){9}
//: {10}(6,124)(6,180)(39,180){11}
//: {12}(210,124)(210,175)(243,175){13}
wire w23;    //: /sn:0 {0}(577,217)(621,217){1}
wire [1:0] w10;    //: /sn:0 {0}(-140,149)(-140,432)(646,432){1}
wire [2:0] w24;    //: /sn:0 {0}(431,193)(381,193)(381,141){1}
//: {2}(383,139)(568,139)(568,193)(621,193){3}
//: {4}(379,139)(260,139)(260,138)(195,138){5}
//: {6}(191,138)(-13,138){7}
//: {8}(-17,138)(-65,138)(-65,-33){9}
//: {10}(-15,140)(-15,193)(39,193){11}
//: {12}(193,140)(193,188)(243,188){13}
wire w31;    //: /sn:0 {0}(243,200)(178,200)(178,60)(100,60)(100,19){1}
wire w1;    //: /sn:0 {0}(-17,217)(39,217){1}
wire [31:0] R1;    //: {0}(281,223)(281,308)(53,308)(53,353){1}
wire [31:0] R3;    //: {0}(687,228)(687,416){1}
wire [1:0] w11;    //: /sn:0 {0}(-27,-33)(-27,-23)(106,-23)(106,-10){1}
wire w2;    //: /sn:0 {0}(243,212)(204,212){1}
wire [31:0] R0;    //: {0}(77,228)(77,299)(41,299)(41,353){1}
wire [31:0] w5;    //: /sn:0 {0}(675,416)(675,372)(497,372)(497,228){1}
wire [31:0] w9;    //: /sn:0 {0}(663,416)(663,387)(309,387)(309,223){1}
//: enddecls

  //: joint g8 (w18) @(6, 122) /w:[ 7 -1 8 10 ]
  //: input g4 (Read2) @(-239,145) /sn:0 /w:[ 0 ]
  //: joint g44 (clr) @(353, -83) /w:[ 3 -1 4 10 ]
  //: input g3 (Write) @(-240,-38) /sn:0 /w:[ 0 ]
  //: joint g16 (clk) @(165, 285) /w:[ 5 6 8 -1 ]
  //: joint g47 (clr) @(541, -83) /w:[ 1 -1 2 12 ]
  //: input g17 (Read1) @(-239,96) /sn:0 /w:[ 0 ]
  //: joint g26 (w19) @(229, 106) /w:[ 5 -1 6 12 ]
  //: output g2 (Data2) @(668,482) /sn:0 /R:3 /w:[ 0 ]
  tran g23(.Z(w24), .I(Write[2:0]));   //: @(-65,-39) /sn:0 /R:1 /w:[ 9 1 2 ] /ss:1
  tran g30(.Z(w10), .I(Read2[4:3]));   //: @(-140,143) /sn:0 /R:1 /w:[ 0 1 2 ] /ss:1
  //: output g1 (Data1) @(59,462) /sn:0 /R:3 /w:[ 1 ]
  //: joint g39 (RegWrite) @(372, 263) /w:[ 6 8 5 -1 ]
  Regs8x32 g24 (.DIN(WriteData), .SD(w24), .SA(w19), .SB(w18), .RegWr(w31), .clk(w2), .clr(clr), .AOUT(R1), .BOUT(w9));   //: @(244, 153) /sz:(98, 69) /sn:0 /p:[ Ti0>11 Li0>13 Li1>13 Li2>13 Li3>0 Li4>0 Ri0>11 Bo0<0 Bo1<1 ]
  Regs8x32 g29 (.DIN(WriteData), .SD(w24), .SA(w19), .SB(w18), .RegWr(w4), .clk(w22), .clr(clr), .AOUT(R2), .BOUT(w5));   //: @(432, 158) /sz:(98, 69) /sn:0 /p:[ Ti0>13 Li0>0 Li1>0 Li2>0 Li3>1 Li4>1 Ri0>13 Bo0<1 Bo1<1 ]
  //: comment g51 /dolink:0 /link:"" @(395,229) /sn:0
  //: /line:"Regs 16-23"
  //: /end
  tran g18(.Z(w19), .I(Read1[2:0]));   //: @(-95,93) /sn:0 /R:1 /w:[ 9 3 4 ] /ss:1
  //: supply1 g10 (w21) @(68,-11) /sn:0 /w:[ 1 ]
  //: joint g25 (w18) @(210, 122) /w:[ 5 -1 6 12 ]
  //: comment g49 /dolink:0 /link:"" @(210,225) /sn:0
  //: /line:"Regs 8-15"
  //: /end
  //: comment g50 /dolink:0 /link:"" @(585,229) /sn:0
  //: /line:"Regs 24-31"
  //: /end
  Regs8x32 g6 (.DIN(WriteData), .SD(w24), .SA(w19), .SB(w18), .RegWr(w16), .clk(w1), .clr(clr), .AOUT(R0), .BOUT(w0));   //: @(40, 158) /sz:(98, 69) /sn:0 /p:[ Ti0>9 Li0>11 Li1>11 Li2>11 Li3>0 Li4>1 Ri0>9 Bo0<0 Bo1<1 ]
  //: joint g7 (w19) @(23, 106) /w:[ 7 -1 8 10 ]
  demux g9 (.I(w11), .E(w21), .Z0(w16), .Z1(w31), .Z2(w4), .Z3(w20));   //: @(106,3) /sn:0 /w:[ 1 0 1 1 0 0 ]
  and g35 (.I0(clk), .I1(RegWrite), .Z(w22));   //: @(394,217) /sn:0 /delay:" 1" /w:[ 3 9 0 ]
  tran g31(.Z(w6), .I(Read1[4:3]));   //: @(-123,93) /sn:0 /R:1 /w:[ 1 1 2 ] /ss:1
  tran g22(.Z(w18), .I(Read2[2:0]));   //: @(-93,142) /sn:0 /R:1 /w:[ 9 3 4 ] /ss:0
  and g36 (.I0(clk), .I1(RegWrite), .Z(w23));   //: @(567,217) /sn:0 /delay:" 1" /w:[ 0 7 0 ]
  //: joint g41 (w19) @(419, 107) /w:[ 2 -1 4 1 ]
  //: joint g45 (WriteData) @(479, 75) /w:[ 1 -1 2 12 ]
  and g33 (.I0(clk), .I1(RegWrite), .Z(w1));   //: @(-27,217) /sn:0 /delay:" 1" /w:[ 11 13 0 ]
  //: input g42 (clr) @(-237,-92) /sn:0 /w:[ 7 ]
  //: joint g40 (w18) @(402, 123) /w:[ 2 -1 4 1 ]
  //: input g12 (clk) @(-239,285) /sn:0 /w:[ 13 ]
  and g34 (.I0(clk), .I1(RegWrite), .Z(w2));   //: @(194,212) /sn:0 /delay:" 1" /w:[ 7 11 1 ]
  //: joint g28 (w24) @(381, 139) /w:[ 2 -1 4 1 ]
  Regs8x32 g46 (.DIN(WriteData), .SD(w24), .SA(w19), .SB(w18), .RegWr(w20), .clk(w23), .clr(clr), .AOUT(w3), .BOUT(R3));   //: @(622, 158) /sz:(98, 69) /sn:0 /p:[ Ti0>0 Li0>3 Li1>3 Li2>3 Li3>1 Li4>1 Ri0>0 Bo0<1 Bo1<0 ]
  //: joint g11 (w24) @(-15, 138) /w:[ 7 -1 8 10 ]
  mux g14 (.I0(R0), .I1(R1), .I2(R2), .I3(w3), .S(w6), .Z(Data1));   //: @(59,369) /sn:0 /w:[ 1 1 0 0 0 0 ] /ss:0 /do:0
  tran g5(.Z(w11), .I(Write[4:3]));   //: @(-27,-39) /sn:0 /R:1 /w:[ 0 3 4 ] /ss:1
  //: joint g19 (clk) @(-58, 285) /w:[ 9 10 12 -1 ]
  //: joint g21 (w24) @(193, 138) /w:[ 5 -1 6 12 ]
  //: input g32 (RegWrite) @(-239,263) /sn:0 /w:[ 0 ]
  //: joint g20 (WriteData) @(87, 75) /w:[ 5 -1 6 8 ]
  //: joint g38 (RegWrite) @(173, 263) /w:[ 4 10 3 -1 ]
  //: joint g15 (clk) @(362, 285) /w:[ 1 2 4 -1 ]
  //: joint g43 (clr) @(148, -83) /w:[ 5 -1 6 8 ]
  //: input g0 (WriteData) @(-239,73) /sn:0 /w:[ 7 ]
  //: joint g27 (WriteData) @(290, 75) /w:[ 3 -1 4 10 ]
  //: comment g48 /dolink:0 /link:"" @(11,228) /sn:0
  //: /line:"Regs 0-7"
  //: /end
  //: joint g37 (RegWrite) @(-69, 263) /w:[ 2 12 1 -1 ]
  mux g13 (.I0(w0), .I1(w9), .I2(w5), .I3(R3), .S(w10), .Z(Data2));   //: @(669,432) /sn:0 /w:[ 0 0 0 1 1 1 ] /ss:0 /do:0

endmodule

module Regs8x32(SB, SA, BOUT, AOUT, clk, clr, RegWr, SD, DIN);
//: interface  /sz:(98, 69) /bd:[ Ti0>DIN[31:0](47/98) Li0>clk(59/69) Li1>RegWr(47/69) Li2>SB[2:0](22/69) Li3>SA[2:0](11/69) Li4>SD[2:0](35/69) Ri0>clr(35/69) Bo0<BOUT[31:0](65/98) Bo1<AOUT[31:0](37/98) ]
input [31:0] DIN;    //: /sn:0 {0}(531,269)(531,318){1}
//: {2}(533,320)(627,320){3}
//: {4}(631,320)(715,320){5}
//: {6}(719,320)(807,320)(807,429){7}
//: {8}(717,322)(717,352){9}
//: {10}(629,322)(629,433){11}
//: {12}(529,320)(435,320){13}
//: {14}(431,320)(342,320){15}
//: {16}(338,320)(264,320){17}
//: {18}(260,320)(181,320)(181,352){19}
//: {20}(262,322)(262,439){21}
//: {22}(340,322)(340,351){23}
//: {24}(433,322)(433,436){25}
//: {26}(531,322)(531,348){27}
output [31:0] BOUT;    //: /sn:0 {0}(516,697)(516,672){1}
input [2:0] SD;    //: /sn:0 {0}(782,138)(852,138)(852,156){1}
supply1 w21;    //: /sn:0 {0}(828,169)(801,169)(801,153){1}
input [2:0] SB;    //: /sn:0 {0}(466,659)(493,659){1}
input RegWr;    //: /sn:0 {0}(48,363)(68,363)(68,378)(82,378){1}
input [2:0] SA;    //: /sn:0 {0}(256,657)(231,657){1}
input clr;    //: /sn:0 /dp:1 {0}(959,337)(1032,337){1}
input clk;    //: /sn:0 {0}(82,383)(68,383)(68,398)(55,398){1}
output [31:0] AOUT;    //: /sn:0 {0}(279,670)(279,702){1}
wire [31:0] w16;    //: /sn:0 {0}(531,369)(531,574)(520,574){1}
//: {2}(516,574)(282,574)(282,641){3}
//: {4}(518,576)(518,587)(519,587)(519,643){5}
wire w7;    //: /sn:0 {0}(472,451)(513,451)(513,405)(848,405)(848,185){1}
wire [31:0] R5;    //: {0}(288,641)(288,586)(525,586){1}
//: {2}(529,586)(629,586)(629,454){3}
//: {4}(527,588)(527,617)(525,617)(525,643){5}
wire w4;    //: /sn:0 {0}(943,337)(906,337){1}
//: {2}(902,337)(767,337){3}
//: {4}(763,337)(588,337){5}
//: {6}(584,337)(390,337){7}
//: {8}(386,337)(231,337)(231,357)(220,357){9}
//: {10}(388,339)(388,356)(379,356){11}
//: {12}(586,339)(586,353)(570,353){13}
//: {14}(765,339)(765,357)(756,357){15}
//: {16}(904,339)(904,417)(865,417){17}
//: {18}(861,417)(675,417){19}
//: {20}(671,417)(489,417){21}
//: {22}(485,417)(302,417)(302,444)(301,444){23}
//: {24}(487,419)(487,441)(472,441){25}
//: {26}(673,419)(673,438)(668,438){27}
//: {28}(863,419)(863,434)(846,434){29}
wire [31:0] R2;    //: {0}(262,641)(262,537){1}
//: {2}(264,535)(499,535)(499,643){3}
//: {4}(262,533)(262,460){5}
wire w0;    //: /sn:0 {0}(770,439)(764,439)(764,481)(579,481){1}
//: {2}(577,479)(577,443)(592,443){3}
//: {4}(575,481)(390,481){5}
//: {6}(388,479)(388,446)(396,446){7}
//: {8}(386,481)(214,481){9}
//: {10}(212,479)(212,449)(225,449){11}
//: {12}(210,481)(125,481)(125,383){13}
//: {14}(127,381)(291,381){15}
//: {16}(295,381)(477,381){17}
//: {18}(481,381)(660,381)(660,362)(680,362){19}
//: {20}(479,379)(479,358)(494,358){21}
//: {22}(293,379)(293,361)(303,361){23}
//: {24}(125,379)(125,362)(144,362){25}
//: {26}(123,381)(103,381){27}
wire w3;    //: /sn:0 {0}(835,185)(835,397)(330,397)(330,454)(301,454){1}
wire [31:0] R7;    //: {0}(807,450)(807,609)(541,609){1}
//: {2}(537,609)(302,609)(302,641){3}
//: {4}(539,611)(539,643){5}
wire w12;    //: /sn:0 {0}(756,367)(787,367)(787,258)(868,258)(868,185){1}
wire w10;    //: /sn:0 {0}(846,444)(875,444)(875,185){1}
wire [31:0] R4;    //: {0}(340,372)(340,545){1}
//: {2}(342,547)(505,547)(505,643){3}
//: {4}(338,547)(268,547)(268,641){5}
wire [31:0] R3;    //: {0}(512,643)(512,559)(435,559){1}
//: {2}(433,557)(433,457){3}
//: {4}(431,559)(275,559)(275,641){5}
wire w8;    //: /sn:0 {0}(220,367)(249,367)(249,213)(828,213)(828,185){1}
wire Z5;    //: /sn:0 {0}(861,185)(861,413)(700,413)(700,448)(668,448){1}
wire w14;    //: /sn:0 {0}(379,366)(414,366)(414,229)(841,229)(841,185){1}
wire [31:0] R0;    //: {0}(492,643)(492,523)(257,523){1}
//: {2}(253,523)(181,523)(181,373){3}
//: {4}(255,525)(255,641){5}
wire w15;    //: /sn:0 {0}(570,363)(608,363)(608,244)(855,244)(855,185){1}
wire [31:0] R10;    //: /sn:0 {0}(295,641)(295,600)(530,600){1}
//: {2}(534,600)(717,600)(717,373){3}
//: {4}(532,602)(532,643){5}
//: enddecls

  //: joint g8 (w16) @(518, 574) /w:[ 1 -1 2 4 ]
  //: input g4 (SB) @(464,659) /sn:0 /w:[ 0 ]
  //: input g3 (SA) @(229,657) /sn:0 /w:[ 1 ]
  //: joint g16 (R3) @(433, 559) /w:[ 1 2 4 -1 ]
  //: joint g17 (R4) @(340, 547) /w:[ 2 1 4 -1 ]
  //: joint g26 (DIN) @(340, 320) /w:[ 15 -1 16 22 ]
  register R5 (.Q(R5), .D(DIN), .EN(Z5), .CLR(w4), .CK(!w0));   //: @(629,443) /w:[ 3 11 1 27 3 ]
  //: output g2 (BOUT) @(516,694) /sn:0 /R:3 /w:[ 0 ]
  //: joint g23 (w4) @(765, 337) /w:[ 3 -1 4 14 ]
  //: joint g30 (w0) @(212, 481) /w:[ 9 10 12 -1 ]
  //: output g1 (AOUT) @(279,699) /sn:0 /R:3 /w:[ 1 ]
  //: joint g39 (DIN) @(262, 320) /w:[ 17 -1 18 20 ]
  //: joint g24 (DIN) @(531, 320) /w:[ 2 1 12 26 ]
  //: joint g29 (w0) @(388, 481) /w:[ 5 6 8 -1 ]
  register R2 (.Q(R4), .D(DIN), .EN(w14), .CLR(w4), .CK(!w0));   //: @(340,361) /w:[ 0 23 0 11 23 ]
  register R7 (.Q(R7), .D(DIN), .EN(w10), .CLR(w4), .CK(!w0));   //: @(807,439) /w:[ 0 7 0 29 0 ]
  //: joint g18 (R2) @(262, 535) /w:[ 2 4 -1 1 ]
  //: supply1 g10 (w21) @(812,153) /sn:0 /w:[ 1 ]
  not g25 (.I(clr), .Z(w4));   //: @(953,337) /sn:0 /R:2 /w:[ 0 0 ]
  //: joint g6 (R7) @(539, 609) /w:[ 1 -1 2 4 ]
  register R6 (.Q(R10), .D(DIN), .EN(w12), .CLR(w4), .CK(!w0));   //: @(717,362) /w:[ 3 9 0 15 19 ]
  //: joint g7 (R10) @(532, 600) /w:[ 2 -1 1 4 ]
  register R4 (.Q(w16), .D(DIN), .EN(w15), .CLR(w4), .CK(!w0));   //: @(531,358) /w:[ 0 27 0 13 21 ]
  demux g9 (.I(SD), .E(w21), .Z0(!w8), .Z1(!w3), .Z2(!w14), .Z3(!w7), .Z4(!w15), .Z5(!Z5), .Z6(!w12), .Z7(!w10));   //: @(852,169) /sn:0 /w:[ 1 0 1 0 1 1 1 0 1 1 ]
  and g35 (.I0(RegWr), .I1(clk), .Z(w0));   //: @(93,381) /sn:0 /delay:" 1" /w:[ 1 0 27 ]
  //: joint g31 (w4) @(863, 417) /w:[ 17 -1 18 28 ]
  //: joint g22 (w4) @(586, 337) /w:[ 5 -1 6 12 ]
  register R3 (.Q(R3), .D(DIN), .EN(w7), .CLR(w4), .CK(!w0));   //: @(433,446) /w:[ 3 25 0 25 7 ]
  register R1 (.Q(R2), .D(DIN), .EN(w3), .CLR(w4), .CK(!w0));   //: @(262,449) /w:[ 5 21 1 23 11 ]
  //: joint g36 (w4) @(904, 337) /w:[ 1 -1 2 16 ]
  //: joint g41 (DIN) @(717, 320) /w:[ 6 -1 5 8 ]
  //: joint g33 (w4) @(673, 417) /w:[ 19 -1 20 26 ]
  //: joint g42 (DIN) @(629, 320) /w:[ 4 -1 3 10 ]
  //: joint g40 (DIN) @(433, 320) /w:[ 13 -1 14 24 ]
  //: joint g12 (w0) @(479, 381) /w:[ 18 20 17 -1 ]
  //: input g34 (clk) @(53,398) /sn:0 /w:[ 1 ]
  //: input g28 (clr) @(1034,337) /sn:0 /R:2 /w:[ 1 ]
  //: joint g11 (w0) @(293, 381) /w:[ 16 22 15 -1 ]
  //: input g5 (RegWr) @(46,363) /sn:0 /w:[ 0 ]
  mux g14 (.I0(R0), .I1(R2), .I2(R4), .I3(R3), .I4(w16), .I5(R5), .I6(R10), .I7(R7), .S(SA), .Z(AOUT));   //: @(279,657) /sn:0 /w:[ 5 0 5 5 3 0 0 3 0 0 ] /ss:0 /do:0
  //: joint g19 (R0) @(255, 523) /w:[ 1 -1 2 4 ]
  //: joint g21 (w4) @(388, 337) /w:[ 7 -1 8 10 ]
  //: joint g32 (w4) @(487, 417) /w:[ 21 -1 22 24 ]
  //: input g20 (SD) @(780,138) /sn:0 /w:[ 0 ]
  register R0 (.Q(R0), .D(DIN), .EN(w8), .CLR(w4), .CK(!w0));   //: @(181,362) /w:[ 3 19 0 9 25 ]
  //: joint g38 (w0) @(577, 481) /w:[ 1 2 4 -1 ]
  //: joint g15 (R5) @(527, 586) /w:[ 2 -1 1 4 ]
  //: input g0 (DIN) @(531,267) /sn:0 /R:3 /w:[ 0 ]
  //: joint g27 (w0) @(125, 381) /w:[ 14 24 26 13 ]
  mux g13 (.I0(R0), .I1(R2), .I2(R4), .I3(R3), .I4(w16), .I5(R5), .I6(R10), .I7(R7), .S(SB), .Z(BOUT));   //: @(516,659) /sn:0 /w:[ 0 3 3 0 5 5 5 5 1 1 ] /ss:0 /do:0

endmodule

module main;    //: root_module
wire w6;    //: /sn:0 {0}(658,340)(658,350){1}
wire w16;    //: /sn:0 /dp:1 {0}(1145,113)(1145,125)(1178,125)(1178,151)(1168,151){1}
wire [31:0] w13;    //: /sn:0 {0}(1307,266)(1018,266){1}
wire [31:0] w7;    //: /sn:0 {0}(766,204)(912,204)(912,230)(922,230){1}
wire [31:0] w4;    //: /sn:0 {0}(617,305)(565,305)(565,540){1}
wire [5:0] w25;    //: /sn:0 {0}(853,68)(853,-19)(876,-19){1}
wire [4:0] w3;    //: /sn:0 {0}(617,265)(504,265){1}
wire [31:0] w22;    //: /sn:0 /dp:1 {0}(1263,69)(1237,69)(1237,20)(1098,20)(1098,71){1}
//: {2}(1100,73)(1131,73){3}
//: {4}(1096,73)(853,73){5}
//: {6}(852,73)(711,73)(711,37){7}
wire w20;    //: /sn:0 {0}(1018,232)(1028,232){1}
wire [31:0] w12;    //: /sn:0 /dp:2 {0}(500,494)(500,449){1}
//: {2}(500,448)(500,265){3}
//: {4}(500,264)(500,229){5}
//: {6}(500,228)(500,189){7}
//: {8}(500,188)(500,-9){9}
//: {10}(500,-10)(500,-57){11}
wire [31:0] w19;    //: /sn:0 /dp:1 {0}(1576,69)(1388,69){1}
wire [3:0] w18;    //: /sn:0 /dp:1 {0}(968,143)(968,199){1}
wire w23;    //: /sn:0 /dp:1 {0}(1279,102)(1279,114)(1280,114)(1280,125){1}
wire [31:0] w10;    //: /sn:0 {0}(1131,105)(1101,105)(1101,448)(828,448){1}
wire [31:0] w24;    //: /sn:0 /dp:1 {0}(1292,79)(1299,79)(1299,79)(1359,79){1}
wire w21;    //: /sn:0 {0}(666,114)(684,114)(684,156){1}
wire [4:0] w1;    //: /sn:0 {0}(617,189)(504,189){1}
wire [31:0] w8;    //: /sn:0 {0}(766,296)(912,296)(912,270)(922,270){1}
wire [31:0] w27;    //: /sn:0 {0}(1160,89)(1263,89){1}
wire [31:0] w28;    //: /sn:0 /dp:1 {0}(882,-14)(1330,-14)(1330,59)(1359,59){1}
wire w14;    //: /sn:0 {0}(23334,9092)(23334,9102){1}
wire w11;    //: /sn:0 {0}(1157,50)(1157,57)(1145,57)(1145,65){1}
wire [4:0] w2;    //: /sn:0 {0}(617,229)(504,229){1}
wire [25:0] w15;    //: /sn:0 {0}(504,-9)(876,-9){1}
wire w5;    //: /sn:0 {0}(726,340)(726,350){1}
wire w26;    //: /sn:0 /dp:1 {0}(1375,92)(1375,116){1}
wire [15:0] w9;    //: /sn:0 {0}(619,449)(504,449){1}
//: enddecls

  ALU g8 (.ALU_OP(w18), .A(w7), .B(w8), .Zero(w20), .Result(w13));   //: @(923, 200) /sz:(94, 87) /sn:0 /p:[ Ti0>1 Li0>1 Li1>1 Ro0<0 Ro1<1 ]
  tran g4(.Z(w3), .I(w12[15:11]));   //: @(498,265) /sn:0 /R:2 /w:[ 1 3 4 ] /ss:1
  tran g3(.Z(w9), .I(w12[15:0]));   //: @(498,449) /sn:0 /R:2 /w:[ 1 1 2 ] /ss:1
  //: dip g16 (w4) @(565,551) /sn:0 /R:2 /w:[ 1 ] /st:0
  concat g17 (.I0(w15), .I1(w25), .Z(w28));   //: @(881,-14) /sn:0 /w:[ 1 1 0 ] /dr:0
  //: dip g26 (w18) @(968,133) /sn:0 /w:[ 0 ] /st:0
  //: dip g2 (w12) @(500,-67) /sn:0 /w:[ 11 ] /st:0
  //: dip g23 (w22) @(711,27) /sn:0 /w:[ 7 ] /st:0
  SignExtend g1 (.D16b(w9), .D32b(w10));   //: @(620, 412) /sz:(207, 73) /sn:0 /p:[ Li0>0 Ro0<1 ]
  //: comment g24 /dolink:0 /link:"" @(656,46) /sn:0
  //: /line:"PCnext"
  //: /end
  //: switch g18 (w16) @(1151,151) /sn:0 /w:[ 1 ] /st:0
  mux g10 (.I0(w24), .I1(w28), .S(w26), .Z(w19));   //: @(1375,69) /sn:0 /R:1 /w:[ 1 1 0 1 ] /ss:0 /do:0
  led g25 (.I(w19));   //: @(1583,69) /sn:0 /R:3 /w:[ 0 ] /type:2
  tran g6(.Z(w1), .I(w12[25:21]));   //: @(498,189) /sn:0 /R:2 /w:[ 1 7 8 ] /ss:1
  mux g9 (.I0(w22), .I1(w27), .S(w23), .Z(w24));   //: @(1279,79) /sn:0 /R:1 /w:[ 0 1 0 0 ] /ss:0 /do:1
  add g7 (.A(w10), .B(w22), .S(w27), .CI(w11), .CO(w16));   //: @(1147,89) /sn:0 /R:1 /w:[ 0 3 0 1 0 ]
  tran g22(.Z(w15), .I(w12[25:0]));   //: @(498,-9) /sn:0 /R:2 /w:[ 0 9 10 ] /ss:1
  //: switch g12 (w26) @(1375,130) /sn:0 /R:1 /w:[ 1 ] /st:0
  //: switch g28 (w21) @(649,114) /sn:0 /w:[ 0 ] /st:0
  //: joint g11 (w22) @(1098, 73) /w:[ 2 1 4 -1 ]
  //: switch g14 (w23) @(1280,139) /sn:0 /R:1 /w:[ 1 ] /st:0
  tran g5(.Z(w2), .I(w12[20:16]));   //: @(498,229) /sn:0 /R:2 /w:[ 1 5 6 ] /ss:1
  led g19 (.I(w11));   //: @(1157,43) /sn:0 /w:[ 0 ] /type:0
  tran g21(.Z(w25), .I(w22[31:26]));   //: @(853,71) /sn:0 /R:1 /w:[ 0 6 5 ] /ss:0
  led g20 (.I(w13));   //: @(1314,266) /sn:0 /R:3 /w:[ 0 ] /type:2
  //: comment g15 /dolink:0 /link:"" @(1267,159) /sn:0
  //: /line:"PCSrc"
  //: /end
  BRegs32x32 g0 (.clr(w21), .WriteData(w4), .Write(w3), .Read2(w2), .Read1(w1), .RegWrite(w6), .clk(w5), .Data2(w8), .Data1(w7));   //: @(618, 157) /sz:(147, 182) /sn:0 /p:[ Ti0>1 Li0>0 Li1>0 Li2>0 Li3>0 Bi0>0 Bi1>0 Ro0<0 Ro1<0 ]
  //: switch g27 (w14) @(23334,9079) /sn:0 /R:3 /w:[ 0 ] /st:0
  //: comment g13 /dolink:0 /link:"" @(1364,152) /sn:0
  //: /line:"JUMP"
  //: /end

endmodule
