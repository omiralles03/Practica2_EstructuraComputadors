//: version "1.8.7"

module JUMP(Jump, PCSrc, SignExt, PCNext, PCin, Inm26);
//: interface  /sz:(118, 106) /bd:[ Ti0>Jump(82/118) Ti1>Jump(63/118) Li0>PCNext[31:0](54/106) Li1>Inm26[25:0](24/106) Li2>SignExt[31:0](82/106) Li3>SignExtOut[31:0](91/106) Li4>PCNext[31:0](57/106) Li5>lnm26[25:0](27/106) Bi0>PCSrc(74/118) Bi1>PCSrc(90/118) Ro0<PCin[31:0](51/106) Ro1<PCin[31:0](52/106) ]
input PCSrc;    //: /sn:0 {0}(535,343)(535,322){1}
input [31:0] SignExt;    //: /sn:0 {0}(345,325)(417,325){1}
input [25:0] Inm26;    //: /sn:0 {0}(569,181)(602,181)(602,209)(631,209){1}
supply0 w12;    //: /sn:0 /dp:1 {0}(440,184)(440,170)(453,170)(453,173){1}
input [31:0] PCNext;    //: /sn:0 {0}(345,293)(383,293){1}
//: {2}(387,293)(417,293){3}
//: {4}(385,291)(385,224)(426,224){5}
output [31:0] PCin;    //: /sn:0 /dp:1 {0}(727,289)(767,289){1}
supply1 w1;    //: /sn:0 {0}(431,265)(431,285){1}
input Jump;    //: /sn:0 {0}(714,335)(714,312){1}
wire [31:0] w7;    //: /sn:0 /dp:1 {0}(548,299)(698,299){1}
wire [5:0] w4;    //: /sn:0 {0}(489,219)(631,219){1}
wire [31:0] w0;    //: /sn:0 {0}(366,192)(426,192){1}
wire w3;    //: /sn:0 /dp:1 {0}(431,349)(431,333){1}
wire [31:0] w11;    //: /sn:0 {0}(519,289)(485,289)(485,219){1}
//: {2}(485,218)(485,208)(455,208){3}
wire [31:0] w2;    //: /sn:0 /dp:1 {0}(446,309)(519,309){1}
wire [31:0] w5;    //: /sn:0 /dp:1 {0}(637,214)(654,214)(654,279)(698,279){1}
wire w9;    //: /sn:0 {0}(440,232)(440,242){1}
//: enddecls

  mux g8 (.I0(w7), .I1(w5), .S(Jump), .Z(PCin));   //: @(714,289) /sn:0 /R:1 /w:[ 1 1 1 0 ] /ss:0 /do:0
  //: input g4 (Jump) @(714,337) /sn:0 /R:1 /w:[ 0 ]
  tran g16(.Z(w4), .I(w11[31:26]));   //: @(483,219) /sn:0 /R:2 /w:[ 0 1 2 ] /ss:1
  //: input g3 (PCSrc) @(535,345) /sn:0 /R:1 /w:[ 0 ]
  //: comment g17 /dolink:0 /link:"" @(419,145) /sn:0
  //: /line:"PC + 1"
  //: /end
  //: input g2 (SignExt) @(343,325) /sn:0 /w:[ 0 ]
  //: input g1 (PCNext) @(343,293) /sn:0 /w:[ 0 ]
  //: comment g18 /dolink:0 /link:"" @(389,396) /sn:0
  //: /line:"PC + SignExt + 1"
  //: /line:""
  //: /end
  led g10 (.I(w3));   //: @(431,356) /sn:0 /R:2 /w:[ 0 ] /type:2
  add g6 (.A(SignExt), .B(PCNext), .S(w2), .CI(w1), .CO(w3));   //: @(433,309) /sn:0 /R:1 /w:[ 1 3 0 1 1 ]
  //: supply0 g9 (w12) @(453,179) /sn:0 /w:[ 1 ]
  mux g7 (.I0(w11), .I1(w2), .S(PCSrc), .Z(w7));   //: @(535,299) /sn:0 /R:1 /w:[ 0 1 1 0 ] /ss:0 /do:1
  concat g12 (.I0(Inm26), .I1(w4), .Z(w5));   //: @(636,214) /sn:0 /w:[ 1 1 0 ] /dr:1
  //: joint g11 (PCNext) @(385, 293) /w:[ 2 4 1 -1 ]
  add g14 (.A(PCNext), .B(w0), .S(w11), .CI(w12), .CO(w9));   //: @(442,208) /sn:0 /R:1 /w:[ 5 1 3 0 0 ]
  //: output g5 (PCin) @(764,289) /sn:0 /w:[ 1 ]
  //: supply1 g15 (w1) @(442,265) /sn:0 /w:[ 0 ]
  //: input g0 (Inm26) @(567,181) /sn:0 /w:[ 0 ]
  //: dip g13 (w0) @(328,192) /sn:0 /R:1 /w:[ 0 ] /st:1

endmodule

module main;    //: root_module
wire [31:0] w7;    //: /sn:0 /dp:1 {0}(692,315)(748,315){1}
wire w4;    //: /sn:0 {0}(854,216)(854,241){1}
wire w3;    //: /sn:0 {0}(844,417)(844,387){1}
wire [31:0] w1;    //: /sn:0 /dp:1 {0}(691,354)(748,354){1}
wire [25:0] w2;    //: /sn:0 /dp:1 {0}(692,278)(748,278){1}
wire [31:0] w5;    //: /sn:0 {0}(970,312)(900,312){1}
//: enddecls

  JUMP g4 (.Jump(w4), .SignExt(w1), .Inm26(w2), .PCNext(w7), .PCSrc(w3), .PCin(w5));   //: @(749, 242) /sz:(150, 144) /sn:0 /p:[ Ti0>1 Li0>1 Li1>1 Li2>1 Bi0>1 Ro0<1 ]
  //: switch g3 (w3) @(844,431) /sn:0 /R:1 /w:[ 0 ] /st:0
  //: dip g2 (w1) @(653,354) /sn:0 /R:1 /w:[ 0 ] /st:0
  //: dip g1 (w7) @(654,315) /sn:0 /R:1 /w:[ 0 ] /st:-805306368
  led g6 (.I(w5));   //: @(977,312) /sn:0 /R:3 /w:[ 0 ] /type:2
  //: switch g5 (w4) @(854,203) /sn:0 /R:3 /w:[ 0 ] /st:1
  //: dip g0 (w2) @(654,278) /sn:0 /R:1 /w:[ 0 ] /st:44813807

endmodule
