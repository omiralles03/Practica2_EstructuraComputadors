//: version "1.8.7"

module main;    //: root_module
supply0 w7;    //: /sn:0 {0}(663,372)(663,362)(648,362)(648,393)(639,393)(639,403){1}
supply0 w3;    //: /sn:0 {0}(928,270)(928,255)(899,255)(899,283){1}
supply0 w5;    //: /sn:0 {0}(881,564)(881,466){1}
wire w6;    //: /sn:0 /dp:1 {0}(899,359)(899,339)(899,339)(899,331){1}
wire w13;    //: /sn:0 {0}(556,377)(629,377)(629,403){1}
wire [31:0] w4;    //: /sn:0 {0}(1192,479)(1192,439)(898,439){1}
wire [31:0] w0;    //: /sn:0 {0}(885,323)(787,323)(787,349){1}
wire w12;    //: /sn:0 /dp:1 {0}(634,479)(634,541)(582,541){1}
wire [31:0] w8;    //: /sn:0 {0}(644,441)(686,441){1}
//: {2}(690,441)(863,441){3}
//: {4}(688,439)(688,291)(885,291){5}
wire [31:0] w2;    //: /sn:0 /dp:1 {0}(914,307)(976,307)(976,232)(592,232)(592,441)(623,441){1}
//: enddecls

  clock g8 (.Z(w12));   //: @(569,541) /sn:0 /w:[ 1 ] /omega:2000 /phi:0 /duty:50
  //: switch g4 (w13) @(539,377) /sn:0 /w:[ 0 ] /st:0
  register g3 (.Q(w8), .D(w2), .EN(w7), .CLR(w13), .CK(w12));   //: @(634,441) /sn:0 /R:1 /w:[ 0 1 1 1 0 ]
  rom g2 (.A(w8), .D(w4), .OE(w5));   //: @(881,440) /sn:0 /w:[ 3 1 1 ]
  led g1 (.I(w4));   //: @(1192,486) /sn:0 /R:2 /w:[ 0 ] /type:3
  led g10 (.I(w6));   //: @(899,366) /sn:0 /R:2 /w:[ 0 ] /type:0
  //: supply0 g6 (w3) @(928,276) /sn:0 /w:[ 0 ]
  //: joint g9 (w8) @(688, 441) /w:[ 2 4 1 -1 ]
  //: dip g7 (w0) @(787,360) /sn:0 /R:2 /w:[ 1 ] /st:0
  //: supply0 g11 (w7) @(663,378) /sn:0 /w:[ 0 ]
  //: supply0 g5 (w5) @(881,570) /sn:0 /w:[ 0 ]
  add g0 (.A(w0), .B(w8), .S(w2), .CI(w3), .CO(w6));   //: @(901,307) /sn:0 /R:1 /w:[ 0 5 0 1 1 ]

endmodule
