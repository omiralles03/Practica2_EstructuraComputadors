//: version "1.8.7"

module CONTROL(ALUOp, ALUSrc, MemRead, funct, op, RegDst, Jump, MemWrite, nsubm, RegWrite, Branch, MemToReg);
//: interface  /sz:(130, 230) /bd:[ Li0>op[5:0](154/230) Li1>funct[5:0](187/230) Ro0<RegWrite(215/230) Ro1<ALUSrc(174/230) Ro2<ALUOp[3:0](137/230) Ro3<MemToReg(113/230) Ro4<MemRead(89/230) Ro5<Branch(66/230) Ro6<Jump(43/230) Ro7<RegDst(23/230) Ro8<MemWrite(158/230) Ro9<nsubm(195/230) ]
output Branch;    //: /sn:0 /dp:15 {0}(1075,393)(936,393){1}
//: {2}(934,391)(934,331){3}
//: {4}(936,329)(1023,329){5}
//: {6}(934,327)(934,285)(1023,285){7}
//: {8}(934,395)(934,476){9}
//: {10}(932,478)(923,478)(923,465){11}
//: {12}(934,480)(934,512)(419,512)(419,371){13}
//: {14}(421,369)(651,369){15}
//: {16}(419,367)(419,285){17}
//: {18}(419,281)(419,254){19}
//: {20}(417,283)(390,283)(390,275){21}
supply0 w3;    //: /sn:0 {0}(1150,376)(1129,376)(1129,393){1}
output ALUSrc;    //: /sn:0 {0}(652,472)(633,472){1}
output MemWrite;    //: /sn:0 {0}(652,447)(353,447){1}
//: {2}(351,445)(351,287){3}
//: {4}(351,283)(351,256){5}
//: {6}(349,285)(335,285)(335,277){7}
//: {8}(351,449)(351,465)(612,465){9}
output RegDst;    //: /sn:0 {0}(1023,334)(959,334){1}
//: {2}(957,332)(957,290)(1023,290){3}
//: {4}(957,336)(957,356){5}
//: {6}(959,358)(1071,358){7}
//: {8}(957,360)(957,410){9}
//: {10}(959,412)(1026,412){11}
//: {12}(957,414)(957,477){13}
//: {14}(959,479)(974,479)(974,471){15}
//: {16}(957,481)(957,520)(211,520)(211,498){17}
//: {18}(213,496)(611,496){19}
//: {20}(211,494)(211,298){21}
//: {22}(213,296)(431,296)(431,318)(651,318){23}
//: {24}(211,294)(211,254){25}
//: {26}(209,296)(188,296)(188,272){27}
output RegWrite;    //: /sn:0 /dp:1 {0}(632,496)(653,496){1}
output [3:0] ALUOp;    //: /sn:0 {0}(1156,361)(1168,361){1}
//: {2}(1172,361)(1191,361){3}
//: {4}(1170,363)(1170,392){5}
output MemRead;    //: /sn:0 /dp:1 {0}(636,395)(651,395){1}
input [5:0] funct;    //: /sn:0 {0}(911,468)(898,468){1}
//: {2}(897,468)(880,468){3}
//: {4}(879,468)(860,468){5}
//: {6}(859,468)(840,468){7}
//: {8}(839,468)(826,468){9}
//: {10}(824,466)(824,417)(818,417){11}
//: {12}(822,468)(809,468){13}
output nsubm;    //: /sn:0 {0}(615,392)(591,392){1}
//: {2}(589,390)(589,298){3}
//: {4}(591,296)(654,296){5}
//: {6}(589,294)(589,254){7}
//: {8}(589,394)(589,480)(612,480){9}
output MemToReg;    //: /sn:0 /dp:1 {0}(615,397)(283,397){1}
//: {2}(281,395)(281,289){3}
//: {4}(281,285)(281,256){5}
//: {6}(279,287)(267,287)(267,276){7}
//: {8}(281,399)(281,425){9}
//: {10}(283,427)(651,427){11}
//: {12}(281,429)(281,468){13}
//: {14}(283,470)(612,470){15}
//: {16}(281,472)(281,491)(611,491){17}
input [5:0] op;    //: /sn:0 {0}(122,179)(158,179){1}
output Jump;    //: /sn:0 {0}(652,344)(480,344)(480,286){1}
//: {2}(480,282)(480,254){3}
//: {4}(478,284)(459,284)(459,276){5}
wire w6;    //: /sn:0 {0}(1091,304)(1112,304)(1112,346)(1150,346){1}
wire w7;    //: /sn:0 {0}(546,233)(546,206){1}
//: {2}(548,204)(601,204)(601,233){3}
//: {4}(544,204)(494,204){5}
//: {6}(490,204)(433,204){7}
//: {8}(429,204)(365,204){9}
//: {10}(361,204)(295,204){11}
//: {12}(291,204)(225,204){13}
//: {14}(221,204)(164,204){15}
//: {16}(223,206)(223,233){17}
//: {18}(293,206)(293,235){19}
//: {20}(363,206)(363,235){21}
//: {22}(431,206)(431,233){23}
//: {24}(492,206)(492,233){25}
wire w4;    //: /sn:0 {0}(1092,356)(1150,356){1}
wire w22;    //: /sn:0 {0}(586,233)(586,174)(533,174){1}
//: {2}(529,174)(479,174){3}
//: {4}(475,174)(418,174){5}
//: {6}(414,174)(350,174){7}
//: {8}(346,174)(280,174){9}
//: {10}(276,174)(210,174){11}
//: {12}(206,174)(164,174){13}
//: {14}(208,176)(208,233){15}
//: {16}(278,176)(278,235){17}
//: {18}(348,176)(348,235){19}
//: {20}(416,176)(416,233){21}
//: {22}(477,176)(477,233){23}
//: {24}(531,176)(531,233){25}
wire w0;    //: /sn:0 /dp:1 {0}(534,254)(534,281){1}
//: {2}(536,283)(701,283)(701,259)(1060,259)(1060,299)(1070,299){3}
//: {4}(532,283)(507,283)(507,276){5}
//: {6}(534,285)(534,473){7}
//: {8}(536,475)(612,475){9}
//: {10}(534,477)(534,501)(611,501){11}
wire w20;    //: /sn:0 {0}(1096,396)(1112,396)(1112,366)(1150,366){1}
wire w19;    //: /sn:0 {0}(871,379)(871,391)(878,391){1}
//: {2}(880,389)(880,355){3}
//: {4}(882,353)(1071,353){5}
//: {6}(880,351)(880,321){7}
//: {8}(882,319)(1023,319){9}
//: {10}(880,317)(880,280)(1023,280){11}
//: {12}(880,393)(880,463){13}
wire w18;    //: /sn:0 {0}(1047,410)(1059,410)(1059,398)(1075,398){1}
wire w23;    //: /sn:0 {0}(581,233)(581,164)(528,164){1}
//: {2}(524,164)(474,164){3}
//: {4}(470,164)(413,164){5}
//: {6}(409,164)(345,164){7}
//: {8}(341,164)(275,164){9}
//: {10}(271,164)(205,164){11}
//: {12}(201,164)(164,164){13}
//: {14}(203,166)(203,233){15}
//: {16}(273,166)(273,235){17}
//: {18}(343,166)(343,235){19}
//: {20}(411,166)(411,233){21}
//: {22}(472,166)(472,233){23}
//: {24}(526,166)(526,233){25}
wire w10;    //: /sn:0 {0}(1023,275)(860,275)(860,312){1}
//: {2}(862,314)(1023,314){3}
//: {4}(860,316)(860,387){5}
//: {6}(858,389)(850,389)(850,379){7}
//: {8}(860,391)(860,405){9}
//: {10}(862,407)(1026,407){11}
//: {12}(860,409)(860,463){13}
wire w24;    //: /sn:0 {0}(576,233)(576,154)(523,154){1}
//: {2}(519,154)(469,154){3}
//: {4}(465,154)(408,154){5}
//: {6}(404,154)(340,154){7}
//: {8}(336,154)(270,154){9}
//: {10}(266,154)(200,154){11}
//: {12}(196,154)(164,154){13}
//: {14}(198,156)(198,233){15}
//: {16}(268,156)(268,235){17}
//: {18}(338,156)(338,235){19}
//: {20}(406,156)(406,233){21}
//: {22}(467,156)(467,233){23}
//: {24}(521,156)(521,233){25}
wire w21;    //: /sn:0 {0}(591,233)(591,184)(538,184){1}
//: {2}(534,184)(484,184){3}
//: {4}(480,184)(423,184){5}
//: {6}(419,184)(355,184){7}
//: {8}(351,184)(285,184){9}
//: {10}(281,184)(215,184){11}
//: {12}(211,184)(164,184){13}
//: {14}(213,186)(213,233){15}
//: {16}(283,186)(283,235){17}
//: {18}(353,186)(353,235){19}
//: {20}(421,186)(421,233){21}
//: {22}(482,186)(482,233){23}
//: {24}(536,186)(536,233){25}
wire w1;    //: /sn:0 {0}(1023,324)(898,324)(898,463){1}
wire w11;    //: /sn:0 {0}(1044,280)(1054,280)(1054,304)(1070,304){1}
wire w15;    //: /sn:0 {0}(1044,321)(1055,321)(1055,309)(1070,309){1}
wire w5;    //: /sn:0 {0}(541,233)(541,196){1}
//: {2}(543,194)(596,194)(596,233){3}
//: {4}(539,194)(489,194){5}
//: {6}(485,194)(428,194){7}
//: {8}(424,194)(360,194){9}
//: {10}(356,194)(290,194){11}
//: {12}(286,194)(220,194){13}
//: {14}(216,194)(164,194){15}
//: {16}(218,196)(218,233){17}
//: {18}(288,196)(288,235){19}
//: {20}(358,196)(358,235){21}
//: {22}(426,196)(426,233){23}
//: {24}(487,196)(487,233){25}
wire w9;    //: /sn:0 /dp:1 {0}(1023,270)(840,270)(840,307){1}
//: {2}(842,309)(1023,309){3}
//: {4}(840,311)(840,386){5}
//: {6}(838,388)(825,388)(825,381){7}
//: {8}(840,390)(840,463){9}
//: enddecls

  and g4 (.I0(w7), .I1(!w5), .I2(w21), .I3(!w22), .I4(w23), .I5(w24), .Z(MemWrite));   //: @(351,246) /sn:0 /R:3 /w:[ 21 21 19 19 19 19 5 ]
  //: comment g8 /dolink:0 /link:"" @(248,237) /sn:0 /R:3
  //: /line:"lw"
  //: /end
  //: comment g116 /dolink:0 /link:"" @(497,242) /sn:0
  //: /line:"nandi"
  //: /end
  //: joint g17 (w22) @(208, 174) /w:[ 11 -1 12 14 ]
  //: joint g30 (w23) @(203, 164) /w:[ 11 -1 12 14 ]
  //: joint g74 (RegDst) @(957, 412) /w:[ 10 9 -1 12 ]
  led g92 (.I(RegDst));   //: @(188,265) /sn:0 /w:[ 27 ] /type:0
  or g130 (.I0(nsubm), .I1(MemToReg), .Z(MemRead));   //: @(626,395) /sn:0 /w:[ 0 0 0 ]
  concat g1 (.I0(w24), .I1(w23), .I2(w22), .I3(w21), .I4(w5), .I5(w7), .Z(op));   //: @(159,179) /sn:0 /R:2 /w:[ 13 13 13 13 15 15 1 ] /dr:0
  //: joint g77 (Branch) @(934, 393) /w:[ 1 2 -1 8 ]
  //: comment g111 /dolink:0 /link:"" @(1025,418) /sn:0
  //: /line:"sub/slt"
  //: /end
  or g51 (.I0(MemWrite), .I1(MemToReg), .I2(w0), .I3(nsubm), .Z(ALUSrc));   //: @(623,472) /sn:0 /w:[ 9 15 9 9 1 ]
  //: comment g70 /dolink:0 /link:"" @(904,429) /sn:0 /R:2
  //: /line:"op0"
  //: /end
  //: comment g10 /dolink:0 /link:"" @(382,241) /sn:0 /R:3
  //: /line:"beq"
  //: /end
  //: joint g25 (w23) @(472, 164) /w:[ 3 -1 4 22 ]
  tran g65(.Z(w9), .I(funct[0]));   //: @(840,466) /sn:0 /R:1 /w:[ 9 8 7 ] /ss:0
  led g103 (.I(w9));   //: @(825,374) /sn:0 /w:[ 7 ] /type:0
  //: output g64 (ALUOp) @(1188,361) /sn:0 /w:[ 3 ]
  //: joint g72 (RegDst) @(957, 358) /w:[ 6 5 -1 8 ]
  //: output g49 (ALUSrc) @(649,472) /sn:0 /w:[ 0 ]
  and g6 (.I0(!w7), .I1(!w5), .I2(!w21), .I3(!w22), .I4(w23), .I5(!w24), .Z(Jump));   //: @(480,244) /sn:0 /R:3 /w:[ 25 25 23 23 23 23 3 ]
  //: comment g7 /dolink:0 /link:"" @(148,238) /sn:0 /R:3
  //: /line:"Tipus R"
  //: /end
  //: joint g35 (w5) @(288, 194) /w:[ 11 -1 12 18 ]
  //: output g56 (MemRead) @(648,395) /sn:0 /w:[ 1 ]
  //: joint g58 (MemWrite) @(351, 447) /w:[ 1 2 -1 8 ]
  //: joint g124 (w22) @(531, 174) /w:[ 1 -1 2 24 ]
  //: joint g98 (Branch) @(419, 283) /w:[ -1 18 20 17 ]
  //: joint g85 (RegDst) @(957, 334) /w:[ 1 2 -1 4 ]
  concat g67 (.I0(w6), .I1(w4), .I2(w20), .I3(w3), .Z(ALUOp));   //: @(1155,361) /sn:0 /w:[ 1 1 1 0 0 ] /dr:1
  //: joint g126 (w24) @(521, 154) /w:[ 1 -1 2 24 ]
  //: joint g54 (MemToReg) @(281, 397) /w:[ 1 2 -1 8 ]
  //: joint g33 (w7) @(223, 204) /w:[ 13 -1 14 16 ]
  //: joint g40 (w7) @(363, 204) /w:[ 9 -1 10 20 ]
  or g52 (.I0(MemToReg), .I1(RegDst), .I2(w0), .Z(RegWrite));   //: @(622,496) /sn:0 /w:[ 17 19 11 0 ]
  and g81 (.I0(!w9), .I1(w10), .I2(!w19), .I3(w1), .I4(!Branch), .I5(RegDst), .Z(w15));   //: @(1034,321) /sn:0 /w:[ 3 3 9 0 5 0 0 ]
  //: joint g12 (w24) @(198, 154) /w:[ 11 -1 12 14 ]
  //: joint g108 (w19) @(880, 391) /w:[ -1 2 1 12 ]
  //: joint g131 (nsubm) @(589, 392) /w:[ 1 2 -1 8 ]
  //: joint g106 (w10) @(860, 389) /w:[ -1 5 6 8 ]
  //: joint g96 (MemWrite) @(351, 285) /w:[ -1 4 6 3 ]
  nand g114 (.I0(w19), .I1(RegDst), .Z(w4));   //: @(1082,356) /sn:0 /w:[ 5 7 0 ]
  //: joint g19 (w22) @(348, 174) /w:[ 7 -1 8 18 ]
  //: joint g117 (w0) @(534, 475) /w:[ 8 7 -1 10 ]
  //: joint g78 (w19) @(880, 353) /w:[ 4 6 -1 3 ]
  //: joint g125 (w23) @(526, 164) /w:[ 1 -1 2 24 ]
  //: comment g113 /dolink:0 /link:"" @(1018,362) /sn:0
  //: /line:"NOT and/or"
  //: /end
  //: input g63 (funct) @(807,468) /sn:0 /w:[ 13 ]
  led g93 (.I(MemToReg));   //: @(267,269) /sn:0 /w:[ 7 ] /type:0
  //: joint g100 (Jump) @(480, 284) /w:[ -1 2 4 1 ]
  led g105 (.I(w10));   //: @(850,372) /sn:0 /w:[ 7 ] /type:0
  //: input g0 (op) @(120,179) /sn:0 /w:[ 0 ]
  //: joint g38 (w23) @(343, 164) /w:[ 7 -1 8 18 ]
  //: output g43 (RegDst) @(648,318) /sn:0 /w:[ 23 ]
  led g101 (.I(ALUOp));   //: @(1170,399) /sn:0 /R:2 /w:[ 5 ] /type:2
  //: joint g48 (MemToReg) @(281, 427) /w:[ 10 9 -1 12 ]
  //: joint g37 (w23) @(273, 164) /w:[ 9 -1 10 16 ]
  and g80 (.I0(w9), .I1(!w10), .I2(w19), .I3(!Branch), .I4(RegDst), .Z(w11));   //: @(1034,280) /sn:0 /w:[ 0 0 11 7 3 0 ]
  led g95 (.I(MemWrite));   //: @(335,270) /sn:0 /w:[ 7 ] /type:0
  and g120 (.I0(w7), .I1(!w5), .I2(w21), .I3(!w22), .I4(w23), .I5(!w24), .Z(nsubm));   //: @(589,244) /sn:0 /R:3 /w:[ 3 3 0 0 0 0 7 ]
  //: joint g122 (w5) @(541, 194) /w:[ 2 -1 4 1 ]
  and g76 (.I0(w10), .I1(RegDst), .Z(w18));   //: @(1037,410) /sn:0 /w:[ 11 11 0 ]
  //: output g44 (Jump) @(649,344) /sn:0 /w:[ 0 ]
  //: joint g75 (w10) @(860, 407) /w:[ 10 9 -1 12 ]
  and g3 (.I0(w7), .I1(!w5), .I2(!w21), .I3(!w22), .I4(w23), .I5(w24), .Z(MemToReg));   //: @(281,246) /sn:0 /R:3 /w:[ 19 19 17 17 17 17 5 ]
  //: joint g16 (w24) @(467, 154) /w:[ 3 -1 4 22 ]
  //: output g47 (MemWrite) @(649,447) /sn:0 /w:[ 0 ]
  //: joint g26 (w21) @(421, 184) /w:[ 5 -1 6 20 ]
  led g90 (.I(Branch));   //: @(923,458) /sn:0 /w:[ 11 ] /type:0
  led g109 (.I(funct));   //: @(811,417) /sn:0 /R:1 /w:[ 11 ] /type:2
  and g2 (.I0(!w7), .I1(!w5), .I2(!w21), .I3(!w22), .I4(!w23), .I5(!w24), .Z(RegDst));   //: @(211,244) /sn:0 /R:3 /w:[ 17 17 15 15 15 15 25 ]
  //: output g128 (nsubm) @(651,296) /sn:0 /w:[ 5 ]
  //: joint g23 (w7) @(492, 204) /w:[ 5 -1 6 24 ]
  //: joint g91 (Branch) @(934, 478) /w:[ -1 9 10 12 ]
  tran g86(.Z(w1), .I(funct[3]));   //: @(898,466) /sn:0 /R:1 /w:[ 1 2 1 ] /ss:0
  //: joint g24 (w21) @(482, 184) /w:[ 3 -1 4 22 ]
  //: joint g39 (w21) @(353, 184) /w:[ 7 -1 8 18 ]
  //: joint g104 (w9) @(840, 388) /w:[ -1 5 6 8 ]
  //: comment g127 /dolink:0 /link:"" @(550,246) /sn:0
  //: /line:"nsubm"
  //: /end
  //: joint g29 (w23) @(411, 164) /w:[ 5 -1 6 20 ]
  //: frame g60 @(92,47) /sn:0 /wi:629 /ht:506 /tx:"Unitat Control"
  //: joint g110 (funct) @(824, 468) /w:[ 9 10 12 -1 ]
  //: joint g121 (w7) @(546, 204) /w:[ 2 -1 4 1 ]
  //: joint g18 (w22) @(278, 174) /w:[ 9 -1 10 16 ]
  //: joint g82 (w9) @(840, 309) /w:[ 2 1 -1 4 ]
  //: joint g94 (MemToReg) @(281, 287) /w:[ -1 4 6 3 ]
  //: joint g119 (w0) @(534, 283) /w:[ 2 1 4 6 ]
  led g107 (.I(w19));   //: @(871,372) /sn:0 /w:[ 0 ] /type:0
  //: output g50 (RegWrite) @(650,496) /sn:0 /w:[ 1 ]
  //: comment g9 /dolink:0 /link:"" @(318,237) /sn:0 /R:3
  //: /line:"sw"
  //: /end
  tran g68(.Z(w10), .I(funct[1]));   //: @(860,466) /sn:0 /R:1 /w:[ 13 6 5 ] /ss:0
  or g73 (.I0(Branch), .I1(w18), .Z(w20));   //: @(1086,396) /sn:0 /w:[ 0 1 0 ]
  //: joint g22 (w5) @(487, 194) /w:[ 5 -1 6 24 ]
  //: joint g31 (w21) @(213, 184) /w:[ 11 -1 12 14 ]
  //: joint g59 (MemToReg) @(281, 470) /w:[ 14 13 -1 16 ]
  or g71 (.I0(w0), .I1(w11), .I2(w15), .Z(w6));   //: @(1081,304) /sn:0 /w:[ 3 1 1 0 ]
  //: joint g102 (ALUOp) @(1170, 361) /w:[ 2 -1 1 4 ]
  //: frame g87 @(753,231) /sn:0 /wi:510 /ht:308 /tx:"ALU Control"
  //: joint g83 (w10) @(860, 314) /w:[ 2 1 -1 4 ]
  led g99 (.I(Jump));   //: @(459,269) /sn:0 /w:[ 5 ] /type:0
  //: joint g36 (w21) @(283, 184) /w:[ 9 -1 10 16 ]
  //: joint g41 (w5) @(358, 194) /w:[ 9 -1 10 20 ]
  //: output g45 (Branch) @(648,369) /sn:0 /w:[ 15 ]
  //: comment g42 /dolink:0 /link:"" @(791,48) /sn:0 /R:3
  //: /line:"         opcode      func      ALUOp   ALUCtrl"
  //: /line:"add     00 0000     10 0000     10      0010"
  //: /line:"sub     00 0000     10 0010     10      0110"
  //: /line:"and     00 0000     10 0100     10      0000"
  //: /line:"or      00 0000     10 0101     10      0001"
  //: /line:"slt     00 0000     10 1010     10      0111"
  //: /line:""
  //: /line:"lw      10 0011     XX XXXX     00      0010"
  //: /line:"sw      10 1011     XX XXXX     00      0010"
  //: /line:"nandi   10 1100     XX XXXX     00      0011"
  //: /line:"nsubm   10 1010     XX XXXX     00      0010"
  //: /line:""
  //: /line:"beq     00 0100     XX XXXX     01      0110"
  //: /line:"j       00 0010     XX XXXX     XX      XXXX"
  //: /end
  tran g69(.Z(w19), .I(funct[2]));   //: @(880,466) /sn:0 /R:1 /w:[ 13 4 3 ] /ss:0
  //: supply0 g66 (w3) @(1129,399) /sn:0 /w:[ 1 ]
  //: joint g28 (w7) @(431, 204) /w:[ 7 -1 8 22 ]
  //: joint g34 (w7) @(293, 204) /w:[ 11 -1 12 18 ]
  //: output g46 (MemToReg) @(648,427) /sn:0 /w:[ 11 ]
  and g5 (.I0(!w7), .I1(!w5), .I2(!w21), .I3(w22), .I4(!w23), .I5(!w24), .Z(Branch));   //: @(419,244) /sn:0 /R:3 /w:[ 23 23 21 21 21 21 19 ]
  //: comment g11 /dolink:0 /link:"" @(453,243) /sn:0 /R:3
  //: /line:"j"
  //: /end
  //: joint g14 (w24) @(338, 154) /w:[ 7 -1 8 18 ]
  //: joint g84 (w19) @(880, 319) /w:[ 8 10 -1 7 ]
  led g118 (.I(w0));   //: @(507,269) /sn:0 /w:[ 5 ] /type:0
  //: comment g112 /dolink:0 /link:"" @(1083,402) /sn:0
  //: /line:"beq"
  //: /end
  //: joint g21 (w22) @(477, 174) /w:[ 3 -1 4 22 ]
  //: joint g61 (Branch) @(419, 369) /w:[ 14 16 -1 13 ]
  //: joint g123 (w21) @(536, 184) /w:[ 1 -1 2 24 ]
  and g115 (.I0(w7), .I1(!w5), .I2(w21), .I3(w22), .I4(!w23), .I5(!w24), .Z(w0));   //: @(534,244) /sn:0 /R:3 /w:[ 0 0 25 25 25 25 0 ]
  //: joint g79 (Branch) @(934, 329) /w:[ 4 6 -1 3 ]
  //: joint g20 (w22) @(416, 174) /w:[ 5 -1 6 20 ]
  //: joint g32 (w5) @(218, 194) /w:[ 13 -1 14 16 ]
  led g97 (.I(Branch));   //: @(390,268) /sn:0 /w:[ 21 ] /type:0
  //: joint g129 (nsubm) @(589, 296) /w:[ 4 6 -1 3 ]
  //: joint g15 (w24) @(406, 154) /w:[ 5 -1 6 20 ]
  //: joint g89 (RegDst) @(957, 479) /w:[ 14 13 -1 16 ]
  //: joint g27 (w5) @(426, 194) /w:[ 7 -1 8 22 ]
  //: comment g62 /dolink:0 /link:"" @(964,428) /sn:0 /R:2
  //: /line:"op1"
  //: /end
  //: joint g55 (RegDst) @(211, 496) /w:[ 18 20 -1 17 ]
  led g88 (.I(RegDst));   //: @(974,464) /sn:0 /w:[ 15 ] /type:0
  //: joint g13 (w24) @(268, 154) /w:[ 9 -1 10 16 ]
  //: joint g53 (RegDst) @(211, 296) /w:[ 22 24 26 21 ]

endmodule

module main;    //: root_module
wire [5:0] w4;    //: /sn:0 /dp:1 {0}(640,48)(717,48){1}
wire [5:0] w0;    //: /sn:0 /dp:1 {0}(642,15)(717,15){1}
wire w3;    //: /sn:0 {0}(849,19)(955,19){1}
wire w30;    //: /sn:0 {0}(849,-96)(952,-96){1}
wire w29;    //: /sn:0 {0}(849,-73)(952,-73){1}
wire w23;    //: /sn:0 /dp:1 {0}(849,-50)(953,-50){1}
wire w31;    //: /sn:0 {0}(849,-116)(952,-116){1}
wire w8;    //: /sn:0 /dp:1 {0}(849,62)(953,62){1}
wire w27;    //: /sn:0 {0}(849,-26)(954,-26){1}
wire w2;    //: /sn:0 {0}(882,130)(882,146)(797,146)(797,92){1}
wire [3:0] w26;    //: /sn:0 {0}(849,-2)(1001,-2){1}
wire w9;    //: /sn:0 {0}(849,35)(954,35){1}
//: enddecls

  led g26 (.I(w29));   //: @(959,-73) /sn:0 /R:3 /w:[ 1 ] /type:0
  led g2 (.I(w2));   //: @(882,123) /sn:0 /w:[ 0 ] /type:0
  led g30 (.I(w27));   //: @(961,-26) /sn:0 /R:3 /w:[ 1 ] /type:0
  led g23 (.I(w30));   //: @(959,-96) /sn:0 /R:3 /w:[ 1 ] /type:0
  //: dip g1 (w4) @(602,48) /sn:0 /R:1 /w:[ 0 ] /st:50
  led g29 (.I(w23));   //: @(960,-50) /sn:0 /R:3 /w:[ 1 ] /type:0
  led g31 (.I(w3));   //: @(962,19) /sn:0 /R:3 /w:[ 1 ] /type:0
  led g33 (.I(w9));   //: @(961,35) /sn:0 /R:3 /w:[ 1 ] /type:0
  led g81 (.I(w26));   //: @(1008,-2) /sn:0 /R:3 /w:[ 1 ] /type:2
  led g21 (.I(w31));   //: @(959,-116) /sn:0 /R:3 /w:[ 1 ] /type:0
  //: dip g0 (w0) @(604,15) /sn:0 /R:1 /w:[ 0 ] /st:42
  CONTROL g38 (.funct(w4), .op(w0), .nsubm(w2), .MemWrite(w3), .RegDst(w31), .Jump(w30), .Branch(w29), .MemRead(w23), .MemToReg(w27), .ALUOp(w26), .ALUSrc(w9), .RegWrite(w8));   //: @(718, -139) /sz:(130, 230) /sn:0 /p:[ Li0>1 Li1>1 Bo0<1 Ro0<0 Ro1<0 Ro2<0 Ro3<0 Ro4<0 Ro5<0 Ro6<0 Ro7<0 Ro8<0 ]
  led g37 (.I(w8));   //: @(960,62) /sn:0 /R:3 /w:[ 1 ] /type:0

endmodule
