//: version "1.8.7"

module JUMP(Jump, PCSrc, SignExt, PCNext, PCin, Inm26);
//: interface  /sz:(118, 106) /bd:[ Ti0>Jump(82/118) Ti1>Jump(63/118) Li0>PCNext[31:0](54/106) Li1>Inm26[25:0](24/106) Li2>SignExt[31:0](82/106) Li3>SignExtOut[31:0](91/106) Li4>PCNext[31:0](57/106) Li5>lnm26[25:0](27/106) Bi0>PCSrc(74/118) Bi1>PCSrc(90/118) Ro0<PCin[31:0](51/106) Ro1<PCin[31:0](52/106) ]
input PCSrc;    //: /sn:0 {0}(535,343)(535,322){1}
input [31:0] SignExt;    //: /sn:0 {0}(345,325)(417,325){1}
input [25:0] Inm26;    //: /sn:0 {0}(569,181)(602,181)(602,209)(631,209){1}
supply0 w12;    //: /sn:0 /dp:1 {0}(440,184)(440,170)(453,170)(453,173){1}
input [31:0] PCNext;    //: /sn:0 {0}(345,293)(383,293){1}
//: {2}(387,293)(417,293){3}
//: {4}(385,291)(385,224)(426,224){5}
output [31:0] PCin;    //: /sn:0 /dp:1 {0}(727,289)(767,289){1}
supply1 w1;    //: /sn:0 {0}(431,265)(431,285){1}
input Jump;    //: /sn:0 {0}(714,335)(714,312){1}
wire [31:0] w7;    //: /sn:0 /dp:1 {0}(548,299)(698,299){1}
wire [5:0] w4;    //: /sn:0 {0}(489,219)(631,219){1}
wire [31:0] w0;    //: /sn:0 {0}(366,192)(426,192){1}
wire w3;    //: /sn:0 /dp:1 {0}(431,349)(431,333){1}
wire [31:0] w11;    //: /sn:0 {0}(519,289)(485,289)(485,219){1}
//: {2}(485,218)(485,208)(455,208){3}
wire [31:0] w2;    //: /sn:0 /dp:1 {0}(446,309)(519,309){1}
wire [31:0] w5;    //: /sn:0 /dp:1 {0}(637,214)(654,214)(654,279)(698,279){1}
wire w9;    //: /sn:0 {0}(440,232)(440,242){1}
//: enddecls

  mux g8 (.I0(w7), .I1(w5), .S(Jump), .Z(PCin));   //: @(714,289) /sn:0 /R:1 /w:[ 1 1 1 0 ] /ss:0 /do:0
  //: input g4 (Jump) @(714,337) /sn:0 /R:1 /w:[ 0 ]
  tran g16(.Z(w4), .I(w11[31:26]));   //: @(483,219) /sn:0 /R:2 /w:[ 0 1 2 ] /ss:1
  //: input g3 (PCSrc) @(535,345) /sn:0 /R:1 /w:[ 0 ]
  //: comment g17 /dolink:0 /link:"" @(419,145) /sn:0
  //: /line:"PC + 1"
  //: /end
  //: input g2 (SignExt) @(343,325) /sn:0 /w:[ 0 ]
  //: input g1 (PCNext) @(343,293) /sn:0 /w:[ 0 ]
  //: comment g18 /dolink:0 /link:"" @(389,396) /sn:0
  //: /line:"PC + SignExt + 1"
  //: /line:""
  //: /end
  led g10 (.I(w3));   //: @(431,356) /sn:0 /R:2 /w:[ 0 ] /type:2
  add g6 (.A(SignExt), .B(PCNext), .S(w2), .CI(w1), .CO(w3));   //: @(433,309) /sn:0 /R:1 /w:[ 1 3 0 1 1 ]
  //: supply0 g9 (w12) @(453,179) /sn:0 /w:[ 1 ]
  mux g7 (.I0(w11), .I1(w2), .S(PCSrc), .Z(w7));   //: @(535,299) /sn:0 /R:1 /w:[ 0 1 1 0 ] /ss:0 /do:1
  concat g12 (.I0(Inm26), .I1(w4), .Z(w5));   //: @(636,214) /sn:0 /w:[ 1 1 0 ] /dr:1
  //: joint g11 (PCNext) @(385, 293) /w:[ 2 4 1 -1 ]
  add g14 (.A(PCNext), .B(w0), .S(w11), .CI(w12), .CO(w9));   //: @(442,208) /sn:0 /R:1 /w:[ 5 1 3 0 0 ]
  //: output g5 (PCin) @(764,289) /sn:0 /w:[ 1 ]
  //: supply1 g15 (w1) @(442,265) /sn:0 /w:[ 0 ]
  //: input g0 (Inm26) @(567,181) /sn:0 /w:[ 0 ]
  //: dip g13 (w0) @(328,192) /sn:0 /R:1 /w:[ 0 ] /st:1

endmodule

module MEM(WriteData, ReadData, Adress, clk, MemRead, MemWrite);
//: interface  /sz:(100, 101) /bd:[ Ti0>MemWrite(51/100) Li0>Adress[31:0](31/101) Li1>WriteData[31:0](74/101) Bi0>MemRead(51/100) Ri0>clk(73/101) Ro0<ReadData[31:0](29/101) ]
output [31:0] ReadData;    //: /sn:0 {0}(619,312)(619,331){1}
//: {2}(621,333)(652,333){3}
//: {4}(617,333)(604,333){5}
input [31:0] WriteData;    //: /sn:0 {0}(619,254)(619,296){1}
supply0 w0;    //: /sn:0 {0}(580,373)(580,360){1}
input [31:0] Adress;    //: /sn:0 {0}(529,335)(569,335){1}
input MemWrite;    //: /sn:0 /dp:1 {0}(546,285)(516,285)(516,245){1}
input clk;    //: /sn:0 {0}(503,290)(546,290){1}
input MemRead;    //: /sn:0 {0}(594,387)(594,360){1}
wire w3;    //: /sn:0 {0}(567,288)(585,288){1}
//: {2}(589,288)(638,288)(638,304)(624,304){3}
//: {4}(587,290)(587,310){5}
//: enddecls

  bufif1 g4 (.Z(ReadData), .I(WriteData), .E(w3));   //: @(619,302) /sn:0 /R:3 /w:[ 0 1 3 ]
  //: supply0 g8 (w0) @(580,379) /sn:0 /w:[ 0 ]
  //: input g3 (WriteData) @(619,252) /sn:0 /R:3 /w:[ 0 ]
  //: output g2 (ReadData) @(649,333) /sn:0 /w:[ 3 ]
  //: input g1 (Adress) @(527,335) /sn:0 /w:[ 0 ]
  //: joint g6 (ReadData) @(619, 333) /w:[ 2 1 4 -1 ]
  //: input g7 (clk) @(501,290) /sn:0 /w:[ 0 ]
  //: input g9 (MemRead) @(594,389) /sn:0 /R:1 /w:[ 0 ]
  //: joint g12 (w3) @(587, 288) /w:[ 2 -1 1 4 ]
  and g11 (.I0(MemWrite), .I1(clk), .Z(w3));   //: @(557,288) /sn:0 /w:[ 0 1 0 ]
  //: input g5 (MemWrite) @(516,243) /sn:0 /R:3 /w:[ 1 ]
  ram g0 (.A(Adress), .D(ReadData), .WE(!w3), .OE(!MemRead), .CS(w0));   //: @(587,334) /sn:0 /w:[ 1 5 5 1 1 ]

endmodule

module READ(Data1, Read2, clr, clk, RegWrite, Write, Read1, WriteData, Data2, RegDst, SignExtOut, SignExtIn);
//: interface  /sz:(173, 238) /bd:[ Ti0>RegWrite(85/173) Ti1>RegWrite(82/173) Ti2>RegWrite(82/173) Ti3>RegWrite(82/173) Li0>Read1[4:0](29/238) Li1>Read2[4:0](70/238) Li2>Write[4:0](106/238) Li3>WriteData[31:0](174/238) Li4>SignExtIn[15:0](205/238) Li5>RegDst(140/238) Li6>SignExtIn[15:0](203/238) Li7>WriteData[31:0](173/238) Li8>RegDst(142/238) Li9>Write[4:0](107/238) Li10>Read2[4:0](70/238) Li11>Read1[4:0](37/238) Li12>Read1[4:0](37/238) Li13>Read2[4:0](70/238) Li14>Write[4:0](107/238) Li15>RegDst(142/238) Li16>WriteData[31:0](173/238) Li17>SignExtIn[15:0](203/238) Li18>Read1[4:0](37/238) Li19>Read2[4:0](70/238) Li20>Write[4:0](107/238) Li21>RegDst(142/238) Li22>WriteData[31:0](173/238) Li23>SignExtIn[15:0](203/238) Bi0>clk(57/173) Bi1>clr(119/173) Bi2>clr(124/173) Bi3>clk(62/173) Bi4>clk(62/173) Bi5>clr(124/173) Bi6>clk(62/173) Bi7>clr(124/173) Ro0<SignExtOut[31:0](208/238) Ro1<Data2[31:0](140/238) Ro2<Data1[31:0](78/238) Ro3<SignExtOut[31:0](200/238) Ro4<Data2[31:0](130/238) Ro5<Data1[31:0](90/238) Ro6<Data1[31:0](90/238) Ro7<Data2[31:0](130/238) Ro8<SignExtOut[31:0](200/238) Ro9<Data1[31:0](90/238) Ro10<Data2[31:0](130/238) Ro11<SignExtOut[31:0](200/238) ]
output [31:0] Data2;    //: /sn:0 {0}(323,263)(353,263){1}
input [4:0] Write;    //: /sn:0 {0}(69,242)(114,242){1}
input [31:0] WriteData;    //: /sn:0 {0}(73,303)(148,303)(148,277)(174,277){1}
output [31:0] Data1;    //: /sn:0 /dp:1 {0}(323,171)(354,171){1}
output [31:0] SignExtOut;    //: /sn:0 /dp:1 {0}(330,391)(352,391){1}
input RegDst;    //: /sn:0 {0}(74,274)(130,274)(130,255){1}
input RegWrite;    //: /sn:0 {0}(215,333)(215,307){1}
input clr;    //: /sn:0 {0}(241,97)(241,123){1}
input clk;    //: /sn:0 {0}(283,335)(283,307){1}
input [4:0] Read1;    //: /sn:0 {0}(73,156)(174,156){1}
input [4:0] Read2;    //: /sn:0 {0}(71,196)(98,196){1}
//: {2}(102,196)(174,196){3}
//: {4}(100,198)(100,222)(114,222){5}
input [15:0] SignExtIn;    //: /sn:0 {0}(138,392)(180,392){1}
wire [4:0] w6;    //: /sn:0 /dp:1 {0}(143,232)(174,232){1}
//: enddecls

  //: output g4 (Data1) @(351,171) /sn:0 /w:[ 1 ]
  //: input g8 (Read2) @(69,196) /sn:0 /w:[ 0 ]
  //: input g3 (clr) @(241,95) /sn:0 /R:3 /w:[ 0 ]
  //: input g2 (clk) @(283,337) /sn:0 /R:1 /w:[ 0 ]
  //: input g1 (RegWrite) @(215,335) /sn:0 /R:1 /w:[ 0 ]
  //: input g10 (Write) @(67,242) /sn:0 /w:[ 0 ]
  //: input g6 (Read1) @(71,156) /sn:0 /w:[ 0 ]
  mux g7 (.I0(Read2), .I1(Write), .S(RegDst), .Z(w6));   //: @(130,232) /sn:0 /R:1 /w:[ 5 1 1 0 ] /ss:0 /do:1
  //: joint g9 (Read2) @(100, 196) /w:[ 2 -1 1 4 ]
  //: input g12 (WriteData) @(71,303) /sn:0 /w:[ 0 ]
  //: output g5 (Data2) @(350,263) /sn:0 /w:[ 1 ]
  //: input g11 (RegDst) @(72,274) /sn:0 /w:[ 0 ]
  //: output g14 (SignExtOut) @(349,391) /sn:0 /w:[ 1 ]
  BRegs32x32 g0 (.clr(clr), .Read1(Read1), .Read2(Read2), .Write(w6), .WriteData(WriteData), .clk(clk), .RegWrite(RegWrite), .Data1(Data1), .Data2(Data2));   //: @(175, 124) /sz:(147, 182) /sn:0 /p:[ Ti0>1 Li0>1 Li1>3 Li2>1 Li3>1 Bi0>1 Bi1>1 Ro0<0 Ro1<0 ]
  SignExtend g15 (.Inm16(SignExtIn), .Inm32(SignExtOut));   //: @(181, 368) /sz:(148, 40) /sn:0 /p:[ Li0>1 Ro0<0 ]
  //: input g13 (SignExtIn) @(136,392) /sn:0 /w:[ 0 ]

endmodule

module SignExtend(Inm32, Inm16);
//: interface  /sz:(207, 73) /bd:[ Li0>lnm16[15:0](37/73) Li1>Inm16[15:0](43/73) Li2>Inm16[15:0](43/73) Li3>Inm16[15:0](43/73) Ro0<D32b[31:0](36/73) Ro1<Inm32[31:0](41/73) Ro2<Inm32[31:0](41/73) Ro3<Inm32[31:0](41/73) ]
output [31:0] Inm32;    //: /sn:0 {0}(283,267)(339,267){1}
input [15:0] Inm16;    //: /sn:0 {0}(20,272)(105,272){1}
//: {2}(106,272)(277,272){3}
wire w18;    //: /sn:0 {0}(106,267)(106,247){1}
//: {2}(108,245)(175,245){3}
//: {4}(106,243)(106,237){5}
//: {6}(108,235)(175,235){7}
//: {8}(106,233)(106,227){9}
//: {10}(108,225)(175,225){11}
//: {12}(106,223)(106,217){13}
//: {14}(108,215)(175,215){15}
//: {16}(106,213)(106,207){17}
//: {18}(108,205)(175,205){19}
//: {20}(106,203)(106,197){21}
//: {22}(108,195)(175,195){23}
//: {24}(106,193)(106,187){25}
//: {26}(108,185)(175,185){27}
//: {28}(106,183)(106,177){29}
//: {30}(108,175)(175,175){31}
//: {32}(106,173)(106,167){33}
//: {34}(108,165)(175,165){35}
//: {36}(106,163)(106,157){37}
//: {38}(108,155)(175,155){39}
//: {40}(106,153)(106,147){41}
//: {42}(108,145)(175,145){43}
//: {44}(106,143)(106,137){45}
//: {46}(108,135)(175,135){47}
//: {48}(106,133)(106,127){49}
//: {50}(108,125)(175,125){51}
//: {52}(106,123)(106,117){53}
//: {54}(108,115)(175,115){55}
//: {56}(106,113)(106,107){57}
//: {58}(108,105)(175,105){59}
//: {60}(106,103)(106,95)(175,95){61}
wire [15:0] w1;    //: /sn:0 /dp:1 {0}(277,262)(227,262)(227,170)(181,170){1}
//: enddecls

  tran g4(.Z(w18), .I(Inm16[15]));   //: @(106,270) /sn:0 /R:1 /w:[ 0 1 2 ] /ss:0
  //: joint g8 (w18) @(106, 215) /w:[ 14 16 -1 13 ]
  //: joint g3 (w18) @(106, 245) /w:[ 2 4 -1 1 ]
  //: joint g16 (w18) @(106, 135) /w:[ 46 48 -1 45 ]
  //: joint g17 (w18) @(106, 125) /w:[ 50 52 -1 49 ]
  concat g2 (.I0(Inm16), .I1(w1), .Z(Inm32));   //: @(282,267) /sn:0 /w:[ 3 0 0 ] /dr:0
  //: output g1 (Inm32) @(336,267) /sn:0 /w:[ 1 ]
  //: joint g18 (w18) @(106, 115) /w:[ 54 56 -1 53 ]
  //: joint g10 (w18) @(106, 195) /w:[ 22 24 -1 21 ]
  concat g6 (.I0(w18), .I1(w18), .I2(w18), .I3(w18), .I4(w18), .I5(w18), .I6(w18), .I7(w18), .I8(w18), .I9(w18), .I10(w18), .I11(w18), .I12(w18), .I13(w18), .I14(w18), .I15(w18), .Z(w1));   //: @(180,170) /sn:0 /w:[ 3 7 11 15 19 23 27 31 35 39 43 47 51 55 59 61 1 ] /dr:0
  //: joint g7 (w18) @(106, 225) /w:[ 10 12 -1 9 ]
  //: joint g9 (w18) @(106, 205) /w:[ 18 20 -1 17 ]
  //: joint g12 (w18) @(106, 175) /w:[ 30 32 -1 29 ]
  //: joint g5 (w18) @(106, 235) /w:[ 6 8 -1 5 ]
  //: joint g11 (w18) @(106, 185) /w:[ 26 28 -1 25 ]
  //: joint g14 (w18) @(106, 155) /w:[ 38 40 -1 37 ]
  //: joint g19 (w18) @(106, 105) /w:[ 58 60 -1 57 ]
  //: input g0 (Inm16) @(18,272) /sn:0 /w:[ 0 ]
  //: joint g15 (w18) @(106, 145) /w:[ 42 44 -1 41 ]
  //: joint g13 (w18) @(106, 165) /w:[ 34 36 -1 33 ]

endmodule

module CONTROL(ALUOp, ALUSrc, MemRead, funct, op, RegDst, Jump, MemWrite, nsubm, RegWrite, Branch, label, w8, ReadTTY, WriteTTY);
//: interface  /sz:(130, 230) /bd:[ Li0>op[5:0](154/230) Li1>funct[5:0](187/230) Bi0>label[15:0](36/130) Ro0<RegWrite(215/230) Ro1<ALUSrc(174/230) Ro2<ALUOp[3:0](137/230) Ro3<MemToReg(113/230) Ro4<MemRead(89/230) Ro5<Branch(66/230) Ro6<Jump(43/230) Ro7<RegDst(23/230) Ro8<MemWrite(158/230) Ro9<nsubm(195/230) ]
output Branch;    //: /sn:0 /dp:15 {0}(1075,393)(936,393){1}
//: {2}(934,391)(934,331){3}
//: {4}(936,329)(1023,329){5}
//: {6}(934,327)(934,285)(1023,285){7}
//: {8}(934,395)(934,476){9}
//: {10}(932,478)(923,478)(923,465){11}
//: {12}(934,480)(934,512)(419,512)(419,371){13}
//: {14}(421,369)(651,369){15}
//: {16}(419,367)(419,285){17}
//: {18}(419,281)(419,254){19}
//: {20}(417,283)(390,283)(390,275){21}
supply0 w3;    //: /sn:0 {0}(1150,376)(1129,376)(1129,393){1}
input [15:0] label;    //: /sn:0 /dp:1 {0}(377,650)(361,650)(361,628)(311,628){1}
output MemWrite;    //: /sn:0 {0}(512,447)(652,447){1}
output ALUSrc;    //: /sn:0 {0}(652,472)(633,472){1}
output RegDst;    //: /sn:0 {0}(1023,334)(959,334){1}
//: {2}(957,332)(957,290)(1023,290){3}
//: {4}(957,336)(957,356){5}
//: {6}(959,358)(1071,358){7}
//: {8}(957,360)(957,410){9}
//: {10}(959,412)(1026,412){11}
//: {12}(957,414)(957,477){13}
//: {14}(959,479)(974,479)(974,471){15}
//: {16}(957,481)(957,520)(211,520)(211,498){17}
//: {18}(213,496)(611,496){19}
//: {20}(211,494)(211,298){21}
//: {22}(213,296)(431,296)(431,318)(651,318){23}
//: {24}(211,294)(211,254){25}
//: {26}(209,296)(188,296)(188,272){27}
output ReadTTY;    //: /sn:0 {0}(539,570)(620,570){1}
output RegWrite;    //: /sn:0 /dp:1 {0}(632,496)(653,496){1}
output w8;    //: /sn:0 {0}(483,394)(283,394){1}
//: {2}(281,392)(281,289){3}
//: {4}(281,285)(281,256){5}
//: {6}(279,287)(267,287)(267,276){7}
//: {8}(281,396)(281,425){9}
//: {10}(283,427)(651,427){11}
//: {12}(281,429)(281,468){13}
//: {14}(283,470)(612,470){15}
//: {16}(281,472)(281,489){17}
//: {18}(283,491)(611,491){19}
//: {20}(281,493)(281,567)(518,567){21}
output [3:0] ALUOp;    //: /sn:0 {0}(1156,361)(1168,361){1}
//: {2}(1172,361)(1191,361){3}
//: {4}(1170,363)(1170,392){5}
output WriteTTY;    //: /sn:0 {0}(621,596)(540,596){1}
input [5:0] funct;    //: /sn:0 {0}(911,468)(898,468){1}
//: {2}(897,468)(880,468){3}
//: {4}(879,468)(860,468){5}
//: {6}(859,468)(840,468){7}
//: {8}(839,468)(826,468){9}
//: {10}(824,466)(824,417)(818,417){11}
//: {12}(822,468)(809,468){13}
output MemRead;    //: /sn:0 /dp:1 {0}(636,395)(651,395){1}
output nsubm;    //: /sn:0 {0}(615,392)(591,392){1}
//: {2}(589,390)(589,298){3}
//: {4}(591,296)(654,296){5}
//: {6}(589,294)(589,254){7}
//: {8}(589,394)(589,480)(612,480){9}
input [5:0] op;    //: /sn:0 {0}(122,179)(158,179){1}
output Jump;    //: /sn:0 {0}(652,344)(480,344)(480,286){1}
//: {2}(480,282)(480,254){3}
//: {4}(478,284)(459,284)(459,276){5}
wire w13;    //: /sn:0 {0}(398,653)(436,653)(436,600){1}
//: {2}(438,598)(519,598){3}
//: {4}(436,596)(436,574){5}
//: {6}(438,572)(518,572){7}
//: {8}(436,570)(436,451){9}
//: {10}(438,449)(491,449){11}
//: {12}(436,447)(436,399)(483,399){13}
wire w6;    //: /sn:0 {0}(1091,304)(1112,304)(1112,346)(1150,346){1}
wire w7;    //: /sn:0 {0}(546,233)(546,206){1}
//: {2}(548,204)(601,204)(601,233){3}
//: {4}(544,204)(494,204){5}
//: {6}(490,204)(433,204){7}
//: {8}(429,204)(365,204){9}
//: {10}(361,204)(295,204){11}
//: {12}(291,204)(225,204){13}
//: {14}(221,204)(164,204){15}
//: {16}(223,206)(223,233){17}
//: {18}(293,206)(293,235){19}
//: {20}(363,206)(363,235){21}
//: {22}(431,206)(431,233){23}
//: {24}(492,206)(492,233){25}
wire w4;    //: /sn:0 {0}(1092,356)(1150,356){1}
wire w0;    //: /sn:0 /dp:1 {0}(534,254)(534,281){1}
//: {2}(536,283)(701,283)(701,259)(1060,259)(1060,299)(1070,299){3}
//: {4}(532,283)(507,283)(507,276){5}
//: {6}(534,285)(534,473){7}
//: {8}(536,475)(612,475){9}
//: {10}(534,477)(534,501)(611,501){11}
wire w22;    //: /sn:0 {0}(586,233)(586,174)(533,174){1}
//: {2}(529,174)(479,174){3}
//: {4}(475,174)(418,174){5}
//: {6}(414,174)(350,174){7}
//: {8}(346,174)(280,174){9}
//: {10}(276,174)(210,174){11}
//: {12}(206,174)(164,174){13}
//: {14}(208,176)(208,233){15}
//: {16}(278,176)(278,235){17}
//: {18}(348,176)(348,235){19}
//: {20}(416,176)(416,233){21}
//: {22}(477,176)(477,233){23}
//: {24}(531,176)(531,233){25}
wire w20;    //: /sn:0 {0}(1096,396)(1112,396)(1112,366)(1150,366){1}
wire w18;    //: /sn:0 {0}(1047,410)(1059,410)(1059,398)(1075,398){1}
wire w19;    //: /sn:0 {0}(871,379)(871,391)(878,391){1}
//: {2}(880,389)(880,355){3}
//: {4}(882,353)(1071,353){5}
//: {6}(880,351)(880,321){7}
//: {8}(882,319)(1023,319){9}
//: {10}(880,317)(880,280)(1023,280){11}
//: {12}(880,393)(880,463){13}
wire w10;    //: /sn:0 {0}(1023,275)(860,275)(860,312){1}
//: {2}(862,314)(1023,314){3}
//: {4}(860,316)(860,387){5}
//: {6}(858,389)(850,389)(850,379){7}
//: {8}(860,391)(860,405){9}
//: {10}(862,407)(1026,407){11}
//: {12}(860,409)(860,463){13}
wire w23;    //: /sn:0 {0}(581,233)(581,164)(528,164){1}
//: {2}(524,164)(474,164){3}
//: {4}(470,164)(413,164){5}
//: {6}(409,164)(345,164){7}
//: {8}(341,164)(275,164){9}
//: {10}(271,164)(205,164){11}
//: {12}(201,164)(164,164){13}
//: {14}(203,166)(203,233){15}
//: {16}(273,166)(273,235){17}
//: {18}(343,166)(343,235){19}
//: {20}(411,166)(411,233){21}
//: {22}(472,166)(472,233){23}
//: {24}(526,166)(526,233){25}
wire w21;    //: /sn:0 {0}(591,233)(591,184)(538,184){1}
//: {2}(534,184)(484,184){3}
//: {4}(480,184)(423,184){5}
//: {6}(419,184)(355,184){7}
//: {8}(351,184)(285,184){9}
//: {10}(281,184)(215,184){11}
//: {12}(211,184)(164,184){13}
//: {14}(213,186)(213,233){15}
//: {16}(283,186)(283,235){17}
//: {18}(353,186)(353,235){19}
//: {20}(421,186)(421,233){21}
//: {22}(482,186)(482,233){23}
//: {24}(536,186)(536,233){25}
wire w24;    //: /sn:0 {0}(576,233)(576,154)(523,154){1}
//: {2}(519,154)(469,154){3}
//: {4}(465,154)(408,154){5}
//: {6}(404,154)(340,154){7}
//: {8}(336,154)(270,154){9}
//: {10}(266,154)(200,154){11}
//: {12}(196,154)(164,154){13}
//: {14}(198,156)(198,233){15}
//: {16}(268,156)(268,235){17}
//: {18}(338,156)(338,235){19}
//: {20}(406,156)(406,233){21}
//: {22}(467,156)(467,233){23}
//: {24}(521,156)(521,233){25}
wire w1;    //: /sn:0 {0}(1023,324)(898,324)(898,463){1}
wire w17;    //: /sn:0 {0}(612,465)(353,465){1}
//: {2}(351,463)(351,446){3}
//: {4}(353,444)(491,444){5}
//: {6}(351,442)(351,287){7}
//: {8}(351,283)(351,256){9}
//: {10}(349,285)(335,285)(335,277){11}
//: {12}(351,467)(351,593)(519,593){13}
wire [15:0] w2;    //: /sn:0 {0}(324,670)(362,670)(362,655)(377,655){1}
wire w11;    //: /sn:0 {0}(1044,280)(1054,280)(1054,304)(1070,304){1}
wire w15;    //: /sn:0 {0}(1044,321)(1055,321)(1055,309)(1070,309){1}
wire w5;    //: /sn:0 {0}(541,233)(541,196){1}
//: {2}(543,194)(596,194)(596,233){3}
//: {4}(539,194)(489,194){5}
//: {6}(485,194)(428,194){7}
//: {8}(424,194)(360,194){9}
//: {10}(356,194)(290,194){11}
//: {12}(286,194)(220,194){13}
//: {14}(216,194)(164,194){15}
//: {16}(218,196)(218,233){17}
//: {18}(288,196)(288,235){19}
//: {20}(358,196)(358,235){21}
//: {22}(426,196)(426,233){23}
//: {24}(487,196)(487,233){25}
wire MemToReg;    //: /sn:0 /dp:1 {0}(615,397)(504,397){1}
wire w9;    //: /sn:0 /dp:1 {0}(1023,270)(840,270)(840,307){1}
//: {2}(842,309)(1023,309){3}
//: {4}(840,311)(840,386){5}
//: {6}(838,388)(825,388)(825,381){7}
//: {8}(840,390)(840,463){9}
//: enddecls

  and g4 (.I0(w7), .I1(!w5), .I2(w21), .I3(!w22), .I4(w23), .I5(w24), .Z(w17));   //: @(351,246) /sn:0 /R:3 /w:[ 21 21 19 19 19 19 9 ]
  //: comment g8 /dolink:0 /link:"" @(248,237) /sn:0 /R:3
  //: /line:"lw"
  //: /end
  //: comment g116 /dolink:0 /link:"" @(497,242) /sn:0
  //: /line:"nandi"
  //: /end
  //: joint g17 (w22) @(208, 174) /w:[ 11 -1 12 14 ]
  and g137 (.I0(w8), .I1(w13), .Z(ReadTTY));   //: @(529,570) /sn:0 /w:[ 21 7 0 ]
  //: joint g30 (w23) @(203, 164) /w:[ 11 -1 12 14 ]
  //: joint g74 (RegDst) @(957, 412) /w:[ 10 9 -1 12 ]
  led g92 (.I(RegDst));   //: @(188,265) /sn:0 /w:[ 27 ] /type:0
  or g130 (.I0(nsubm), .I1(MemToReg), .Z(MemRead));   //: @(626,395) /sn:0 /w:[ 0 0 0 ]
  concat g1 (.I0(w24), .I1(w23), .I2(w22), .I3(w21), .I4(w5), .I5(w7), .Z(op));   //: @(159,179) /sn:0 /R:2 /w:[ 13 13 13 13 15 15 1 ] /dr:0
  //: joint g77 (Branch) @(934, 393) /w:[ 1 2 -1 8 ]
  //: comment g111 /dolink:0 /link:"" @(1025,418) /sn:0
  //: /line:"sub/slt"
  //: /end
  //: joint g144 (w13) @(436, 598) /w:[ 2 4 -1 1 ]
  or g51 (.I0(w17), .I1(w8), .I2(w0), .I3(nsubm), .Z(ALUSrc));   //: @(623,472) /sn:0 /w:[ 0 15 9 9 1 ]
  //: comment g70 /dolink:0 /link:"" @(904,429) /sn:0 /R:2
  //: /line:"op0"
  //: /end
  //: comment g10 /dolink:0 /link:"" @(382,241) /sn:0 /R:3
  //: /line:"beq"
  //: /end
  //: joint g25 (w23) @(472, 164) /w:[ 3 -1 4 22 ]
  tran g65(.Z(w9), .I(funct[0]));   //: @(840,466) /sn:0 /R:1 /w:[ 9 8 7 ] /ss:0
  led g103 (.I(w9));   //: @(825,374) /sn:0 /w:[ 7 ] /type:0
  //: output g64 (ALUOp) @(1188,361) /sn:0 /w:[ 3 ]
  //: joint g72 (RegDst) @(957, 358) /w:[ 6 5 -1 8 ]
  //: output g49 (ALUSrc) @(649,472) /sn:0 /w:[ 0 ]
  and g142 (.I0(w17), .I1(w13), .Z(WriteTTY));   //: @(530,596) /sn:0 /w:[ 13 3 1 ]
  and g136 (.I0(w8), .I1(!w13), .Z(MemToReg));   //: @(494,397) /sn:0 /w:[ 0 13 1 ]
  and g6 (.I0(!w7), .I1(!w5), .I2(!w21), .I3(!w22), .I4(w23), .I5(!w24), .Z(Jump));   //: @(480,244) /sn:0 /R:3 /w:[ 25 25 23 23 23 23 3 ]
  //: joint g58 (w17) @(351, 444) /w:[ 4 6 -1 3 ]
  //: comment g7 /dolink:0 /link:"" @(148,238) /sn:0 /R:3
  //: /line:"Tipus R"
  //: /end
  //: joint g35 (w5) @(288, 194) /w:[ 11 -1 12 18 ]
  //: output g56 (MemRead) @(648,395) /sn:0 /w:[ 1 ]
  //: joint g124 (w22) @(531, 174) /w:[ 1 -1 2 24 ]
  //: joint g98 (Branch) @(419, 283) /w:[ -1 18 20 17 ]
  //: joint g85 (RegDst) @(957, 334) /w:[ 1 2 -1 4 ]
  concat g67 (.I0(w6), .I1(w4), .I2(w20), .I3(w3), .Z(ALUOp));   //: @(1155,361) /sn:0 /w:[ 1 1 1 0 0 ] /dr:1
  //: joint g126 (w24) @(521, 154) /w:[ 1 -1 2 24 ]
  //: joint g54 (w8) @(281, 394) /w:[ 1 2 -1 8 ]
  //: joint g33 (w7) @(223, 204) /w:[ 13 -1 14 16 ]
  //: joint g40 (w7) @(363, 204) /w:[ 9 -1 10 20 ]
  or g52 (.I0(w8), .I1(RegDst), .I2(w0), .Z(RegWrite));   //: @(622,496) /sn:0 /w:[ 19 19 11 0 ]
  and g81 (.I0(!w9), .I1(w10), .I2(!w19), .I3(w1), .I4(!Branch), .I5(RegDst), .Z(w15));   //: @(1034,321) /sn:0 /w:[ 3 3 9 0 5 0 0 ]
  //: dip g132 (w2) @(286,670) /sn:0 /R:1 /w:[ 0 ] /st:-1
  //: joint g12 (w24) @(198, 154) /w:[ 11 -1 12 14 ]
  //: joint g108 (w19) @(880, 391) /w:[ -1 2 1 12 ]
  //: joint g131 (nsubm) @(589, 392) /w:[ 1 2 -1 8 ]
  //: joint g106 (w10) @(860, 389) /w:[ -1 5 6 8 ]
  //: joint g96 (w17) @(351, 285) /w:[ -1 8 10 7 ]
  nand g114 (.I0(w19), .I1(RegDst), .Z(w4));   //: @(1082,356) /sn:0 /w:[ 5 7 0 ]
  //: joint g19 (w22) @(348, 174) /w:[ 7 -1 8 18 ]
  //: joint g117 (w0) @(534, 475) /w:[ 8 7 -1 10 ]
  //: joint g78 (w19) @(880, 353) /w:[ 4 6 -1 3 ]
  //: joint g125 (w23) @(526, 164) /w:[ 1 -1 2 24 ]
  //: comment g113 /dolink:0 /link:"" @(1018,362) /sn:0
  //: /line:"NOT and/or"
  //: /end
  //: input g63 (funct) @(807,468) /sn:0 /w:[ 13 ]
  led g93 (.I(w8));   //: @(267,269) /sn:0 /w:[ 7 ] /type:0
  //: joint g100 (Jump) @(480, 284) /w:[ -1 2 4 1 ]
  led g105 (.I(w10));   //: @(850,372) /sn:0 /w:[ 7 ] /type:0
  //: input g0 (op) @(120,179) /sn:0 /w:[ 0 ]
  //: joint g38 (w23) @(343, 164) /w:[ 7 -1 8 18 ]
  //: output g43 (RegDst) @(648,318) /sn:0 /w:[ 23 ]
  led g101 (.I(ALUOp));   //: @(1170,399) /sn:0 /R:2 /w:[ 5 ] /type:2
  //: joint g48 (w8) @(281, 427) /w:[ 10 9 -1 12 ]
  //: joint g37 (w23) @(273, 164) /w:[ 9 -1 10 16 ]
  and g80 (.I0(w9), .I1(!w10), .I2(w19), .I3(!Branch), .I4(RegDst), .Z(w11));   //: @(1034,280) /sn:0 /w:[ 0 0 11 7 3 0 ]
  led g95 (.I(w17));   //: @(335,270) /sn:0 /w:[ 11 ] /type:0
  and g120 (.I0(w7), .I1(!w5), .I2(w21), .I3(!w22), .I4(w23), .I5(!w24), .Z(nsubm));   //: @(589,244) /sn:0 /R:3 /w:[ 3 3 0 0 0 0 7 ]
  //: joint g122 (w5) @(541, 194) /w:[ 2 -1 4 1 ]
  and g76 (.I0(w10), .I1(RegDst), .Z(w18));   //: @(1037,410) /sn:0 /w:[ 11 11 0 ]
  //: output g44 (Jump) @(649,344) /sn:0 /w:[ 0 ]
  //: joint g75 (w10) @(860, 407) /w:[ 10 9 -1 12 ]
  and g3 (.I0(w7), .I1(!w5), .I2(!w21), .I3(!w22), .I4(w23), .I5(w24), .Z(w8));   //: @(281,246) /sn:0 /R:3 /w:[ 19 19 17 17 17 17 5 ]
  //: joint g16 (w24) @(467, 154) /w:[ 3 -1 4 22 ]
  //: output g47 (MemWrite) @(649,447) /sn:0 /w:[ 1 ]
  //: joint g143 (w17) @(351, 465) /w:[ 1 2 -1 12 ]
  //: joint g26 (w21) @(421, 184) /w:[ 5 -1 6 20 ]
  led g90 (.I(Branch));   //: @(923,458) /sn:0 /w:[ 11 ] /type:0
  led g109 (.I(funct));   //: @(811,417) /sn:0 /R:1 /w:[ 11 ] /type:2
  and g2 (.I0(!w7), .I1(!w5), .I2(!w21), .I3(!w22), .I4(!w23), .I5(!w24), .Z(RegDst));   //: @(211,244) /sn:0 /R:3 /w:[ 17 17 15 15 15 15 25 ]
  //: output g128 (nsubm) @(651,296) /sn:0 /w:[ 5 ]
  //: joint g23 (w7) @(492, 204) /w:[ 5 -1 6 24 ]
  //: joint g91 (Branch) @(934, 478) /w:[ -1 9 10 12 ]
  //: joint g141 (w13) @(436, 449) /w:[ 10 12 -1 9 ]
  tran g86(.Z(w1), .I(funct[3]));   //: @(898,466) /sn:0 /R:1 /w:[ 1 2 1 ] /ss:0
  //: joint g24 (w21) @(482, 184) /w:[ 3 -1 4 22 ]
  //: joint g39 (w21) @(353, 184) /w:[ 7 -1 8 18 ]
  //: joint g104 (w9) @(840, 388) /w:[ -1 5 6 8 ]
  //: comment g127 /dolink:0 /link:"" @(550,246) /sn:0
  //: /line:"nsubm"
  //: /end
  //: joint g29 (w23) @(411, 164) /w:[ 5 -1 6 20 ]
  //: frame g60 @(92,47) /sn:0 /wi:638 /ht:667 /tx:"Unitat Control"
  //: joint g110 (funct) @(824, 468) /w:[ 9 10 12 -1 ]
  //: joint g121 (w7) @(546, 204) /w:[ 2 -1 4 1 ]
  //: joint g18 (w22) @(278, 174) /w:[ 9 -1 10 16 ]
  //: joint g82 (w9) @(840, 309) /w:[ 2 1 -1 4 ]
  //: joint g94 (w8) @(281, 287) /w:[ -1 4 6 3 ]
  //: joint g119 (w0) @(534, 283) /w:[ 2 1 4 6 ]
  led g107 (.I(w19));   //: @(871,372) /sn:0 /w:[ 0 ] /type:0
  //: output g50 (RegWrite) @(650,496) /sn:0 /w:[ 1 ]
  xnor g133 (.I0(label), .I1(w2), .Z(w13));   //: @(388,653) /sn:0 /w:[ 0 1 0 ]
  //: comment g9 /dolink:0 /link:"" @(318,237) /sn:0 /R:3
  //: /line:"sw"
  //: /end
  tran g68(.Z(w10), .I(funct[1]));   //: @(860,466) /sn:0 /R:1 /w:[ 13 6 5 ] /ss:0
  or g73 (.I0(Branch), .I1(w18), .Z(w20));   //: @(1086,396) /sn:0 /w:[ 0 1 0 ]
  //: joint g22 (w5) @(487, 194) /w:[ 5 -1 6 24 ]
  //: joint g31 (w21) @(213, 184) /w:[ 11 -1 12 14 ]
  //: joint g59 (w8) @(281, 470) /w:[ 14 13 -1 16 ]
  or g71 (.I0(w0), .I1(w11), .I2(w15), .Z(w6));   //: @(1081,304) /sn:0 /w:[ 3 1 1 0 ]
  //: joint g102 (ALUOp) @(1170, 361) /w:[ 2 -1 1 4 ]
  //: frame g87 @(753,231) /sn:0 /wi:510 /ht:308 /tx:"ALU Control"
  //: joint g83 (w10) @(860, 314) /w:[ 2 1 -1 4 ]
  led g99 (.I(Jump));   //: @(459,269) /sn:0 /w:[ 5 ] /type:0
  //: joint g36 (w21) @(283, 184) /w:[ 9 -1 10 16 ]
  //: joint g41 (w5) @(358, 194) /w:[ 9 -1 10 20 ]
  //: output g45 (Branch) @(648,369) /sn:0 /w:[ 15 ]
  //: joint g138 (w13) @(436, 572) /w:[ 6 8 -1 5 ]
  //: comment g42 /dolink:0 /link:"" @(791,48) /sn:0 /R:3
  //: /line:"         opcode      func      ALUOp   ALUCtrl"
  //: /line:"add     00 0000     10 0000     10      0010"
  //: /line:"sub     00 0000     10 0010     10      0110"
  //: /line:"and     00 0000     10 0100     10      0000"
  //: /line:"or      00 0000     10 0101     10      0001"
  //: /line:"slt     00 0000     10 1010     10      0111"
  //: /line:""
  //: /line:"lw      10 0011     XX XXXX     00      0010"
  //: /line:"sw      10 1011     XX XXXX     00      0010"
  //: /line:"nandi   10 1100     XX XXXX     00      0011"
  //: /line:"nsubm   10 1010     XX XXXX     00      0010"
  //: /line:""
  //: /line:"beq     00 0100     XX XXXX     01      0110"
  //: /line:"j       00 0010     XX XXXX     XX      XXXX"
  //: /end
  tran g69(.Z(w19), .I(funct[2]));   //: @(880,466) /sn:0 /R:1 /w:[ 13 4 3 ] /ss:0
  //: supply0 g66 (w3) @(1129,399) /sn:0 /w:[ 1 ]
  //: input g57 (label) @(309,628) /sn:0 /w:[ 1 ]
  //: joint g28 (w7) @(431, 204) /w:[ 7 -1 8 22 ]
  //: joint g34 (w7) @(293, 204) /w:[ 11 -1 12 18 ]
  //: output g46 (w8) @(648,427) /sn:0 /w:[ 11 ]
  and g5 (.I0(!w7), .I1(!w5), .I2(!w21), .I3(w22), .I4(!w23), .I5(!w24), .Z(Branch));   //: @(419,244) /sn:0 /R:3 /w:[ 23 23 21 21 21 21 19 ]
  //: comment g11 /dolink:0 /link:"" @(453,243) /sn:0 /R:3
  //: /line:"j"
  //: /end
  //: joint g14 (w24) @(338, 154) /w:[ 7 -1 8 18 ]
  //: joint g84 (w19) @(880, 319) /w:[ 8 10 -1 7 ]
  led g118 (.I(w0));   //: @(507,269) /sn:0 /w:[ 5 ] /type:0
  //: comment g112 /dolink:0 /link:"" @(1083,402) /sn:0
  //: /line:"beq"
  //: /end
  //: joint g21 (w22) @(477, 174) /w:[ 3 -1 4 22 ]
  //: joint g61 (Branch) @(419, 369) /w:[ 14 16 -1 13 ]
  //: joint g123 (w21) @(536, 184) /w:[ 1 -1 2 24 ]
  and g115 (.I0(w7), .I1(!w5), .I2(w21), .I3(w22), .I4(!w23), .I5(!w24), .Z(w0));   //: @(534,244) /sn:0 /R:3 /w:[ 0 0 25 25 25 25 0 ]
  //: joint g79 (Branch) @(934, 329) /w:[ 4 6 -1 3 ]
  //: joint g20 (w22) @(416, 174) /w:[ 5 -1 6 20 ]
  //: joint g32 (w5) @(218, 194) /w:[ 13 -1 14 16 ]
  //: output g134 (ReadTTY) @(617,570) /sn:0 /w:[ 1 ]
  led g97 (.I(Branch));   //: @(390,268) /sn:0 /w:[ 21 ] /type:0
  //: joint g129 (nsubm) @(589, 296) /w:[ 4 6 -1 3 ]
  //: joint g15 (w24) @(406, 154) /w:[ 5 -1 6 20 ]
  //: joint g89 (RegDst) @(957, 479) /w:[ 14 13 -1 16 ]
  //: joint g27 (w5) @(426, 194) /w:[ 7 -1 8 22 ]
  //: comment g62 /dolink:0 /link:"" @(964,428) /sn:0 /R:2
  //: /line:"op1"
  //: /end
  //: joint g55 (RegDst) @(211, 496) /w:[ 18 20 -1 17 ]
  led g88 (.I(RegDst));   //: @(974,464) /sn:0 /w:[ 15 ] /type:0
  and g140 (.I0(w17), .I1(!w13), .Z(MemWrite));   //: @(502,447) /sn:0 /w:[ 5 11 0 ]
  //: joint g139 (w8) @(281, 491) /w:[ 18 17 -1 20 ]
  //: output g135 (WriteTTY) @(618,596) /sn:0 /w:[ 0 ]
  //: joint g53 (RegDst) @(211, 296) /w:[ 22 24 26 21 ]
  //: joint g13 (w24) @(268, 154) /w:[ 9 -1 10 16 ]

endmodule

module ALU(ALU_OP, Zero, ALU_RES, B, A);
//: interface  /sz:(99, 90) /bd:[ Ti0>ALU_OP[3:0](35/99) Li0>B[31:0](68/90) Li1>A[31:0](20/90) Ro0<ALU_RES[31:0](65/90) Ro1<Zero(22/90) ]
input [31:0] B;    //: /sn:0 {0}(358,122)(358,181){1}
//: {2}(360,183)(446,183){3}
//: {4}(358,185)(358,207){5}
//: {6}(360,209)(447,209){7}
//: {8}(358,211)(358,280){9}
//: {10}(360,282)(445,282){11}
//: {12}(358,284)(358,462)(460,462){13}
output Zero;    //: /sn:0 {0}(799,345)(776,345){1}
supply0 w4;    //: /sn:0 {0}(599,451)(621,451){1}
//: {2}(625,451)(631,451){3}
//: {4}(635,451)(641,451){5}
//: {6}(645,451)(651,451){7}
//: {8}(655,451)(661,451){9}
//: {10}(665,451)(671,451){11}
//: {12}(675,451)(681,451){13}
//: {14}(685,451)(691,451){15}
//: {16}(695,451)(701,451){17}
//: {18}(705,451)(711,451){19}
//: {20}(715,451)(721,451){21}
//: {22}(725,451)(731,451){23}
//: {24}(735,451)(741,451){25}
//: {26}(745,451)(751,451){27}
//: {28}(755,451)(761,451){29}
//: {30}(765,451)(771,451){31}
//: {32}(775,451)(781,451){33}
//: {34}(785,451)(791,451){35}
//: {36}(795,451)(801,451){37}
//: {38}(805,451)(811,451){39}
//: {40}(815,451)(821,451){41}
//: {42}(825,451)(831,451){43}
//: {44}(835,451)(841,451){45}
//: {46}(845,451)(851,451){47}
//: {48}(855,451)(861,451){49}
//: {50}(865,451)(871,451){51}
//: {52}(875,451)(881,451){53}
//: {54}(885,451)(891,451){55}
//: {56}(895,451)(901,451){57}
//: {58}(905,451)(911,451){59}
//: {60}(915,451)(923,451)(923,420){61}
//: {62}(913,449)(913,420){63}
//: {64}(903,449)(903,420){65}
//: {66}(893,449)(893,420){67}
//: {68}(883,449)(883,420){69}
//: {70}(873,449)(873,420){71}
//: {72}(863,449)(863,420){73}
//: {74}(853,449)(853,420){75}
//: {76}(843,449)(843,420){77}
//: {78}(833,449)(833,420){79}
//: {80}(823,449)(823,420){81}
//: {82}(813,449)(813,420){83}
//: {84}(803,449)(803,420){85}
//: {86}(793,449)(793,420){87}
//: {88}(783,449)(783,420){89}
//: {90}(773,449)(773,420){91}
//: {92}(763,449)(763,420){93}
//: {94}(753,449)(753,420){95}
//: {96}(743,449)(743,420){97}
//: {98}(733,449)(733,420){99}
//: {100}(723,449)(723,420){101}
//: {102}(713,449)(713,420){103}
//: {104}(703,449)(703,420){105}
//: {106}(693,449)(693,420){107}
//: {108}(683,449)(683,420){109}
//: {110}(673,449)(673,420){111}
//: {112}(663,449)(663,420){113}
//: {114}(653,449)(653,420){115}
//: {116}(643,449)(643,420){117}
//: {118}(633,449)(633,420){119}
//: {120}(623,449)(623,420){121}
output [31:0] ALU_RES;    //: /sn:0 /dp:1 {0}(716,314)(740,314){1}
//: {2}(744,314)(779,314){3}
//: {4}(742,316)(742,345)(755,345){5}
input [31:0] A;    //: /sn:0 /dp:1 {0}(316,128)(316,176){1}
//: {2}(318,178)(446,178){3}
//: {4}(316,180)(316,202){5}
//: {6}(318,204)(447,204){7}
//: {8}(316,206)(316,248){9}
//: {10}(318,250)(445,250){11}
//: {12}(316,252)(316,430)(460,430){13}
supply1 w1;    //: /sn:0 {0}(474,407)(474,422){1}
input [3:0] ALU_OP;    //: /sn:0 {0}(710,226)(710,250)(703,250){1}
//: {2}(702,250)(697,250){3}
supply0 w5;    //: /sn:0 /dp:1 {0}(459,242)(459,228)(482,228)(482,238){1}
wire w6;    //: /sn:0 /dp:1 {0}(459,305)(459,290){1}
wire [31:0] w13;    //: /sn:0 {0}(614,317)(633,317){1}
//: {2}(637,317)(687,317){3}
//: {4}(635,319)(635,323)(687,323){5}
wire [31:0] w7;    //: /sn:0 /dp:1 {0}(467,181)(664,181)(664,288){1}
//: {2}(666,290)(687,290){3}
//: {4}(664,292)(664,310)(687,310){5}
wire w3;    //: /sn:0 {0}(564,402)(564,465)(933,465)(933,420){1}
wire [2:0] w0;    //: /sn:0 {0}(703,254)(703,291){1}
wire [31:0] w18;    //: /sn:0 /dp:1 {0}(687,337)(650,337)(650,396)(778,396)(778,414){1}
wire [31:0] w17;    //: /sn:0 /dp:3 {0}(489,446)(510,446)(510,398)(563,398){1}
//: {2}(564,398)(635,398)(635,330)(687,330){3}
wire [31:0] w2;    //: /sn:0 {0}(474,266)(634,266)(634,303)(687,303){1}
wire w11;    //: /sn:0 /dp:1 {0}(474,486)(474,470){1}
wire [31:0] w9;    //: /sn:0 /dp:1 {0}(687,297)(649,297)(649,207)(468,207){1}
//: enddecls

  //: input g4 (ALU_OP) @(710,224) /sn:0 /R:3 /w:[ 0 ]
  and g8 (.I0(A), .I1(B), .Z(w7));   //: @(457,181) /sn:0 /w:[ 3 3 0 ]
  //: joint g44 (w4) @(883, 451) /w:[ 54 68 53 -1 ]
  //: supply1 g16 (w1) @(485,407) /sn:0 /w:[ 0 ]
  //: output g3 (Zero) @(796,345) /sn:0 /w:[ 0 ]
  //: joint g47 (w4) @(843, 451) /w:[ 46 76 45 -1 ]
  add g17 (.A(!B), .B(A), .S(w17), .CI(w1), .CO(w11));   //: @(476,446) /sn:0 /R:1 /w:[ 13 13 0 1 1 ]
  led g26 (.I(w6));   //: @(459,312) /sn:0 /R:2 /w:[ 0 ] /type:2
  //: output g2 (ALU_RES) @(776,314) /sn:0 /w:[ 3 ]
  nor g23 (.I0(ALU_RES), .Z(Zero));   //: @(766,345) /sn:0 /w:[ 5 1 ]
  //: joint g30 (w4) @(903, 451) /w:[ 58 64 57 -1 ]
  //: input g1 (B) @(358,120) /sn:0 /R:3 /w:[ 0 ]
  //: joint g24 (ALU_RES) @(742, 314) /w:[ 2 -1 1 4 ]
  //: joint g39 (w4) @(793, 451) /w:[ 36 86 35 -1 ]
  //: joint g29 (w4) @(913, 451) /w:[ 60 62 59 -1 ]
  led g60 (.I(w11));   //: @(474,493) /sn:0 /R:2 /w:[ 0 ] /type:2
  //: joint g51 (w4) @(763, 451) /w:[ 30 92 29 -1 ]
  //: dip g18 (w13) @(576,317) /sn:0 /R:1 /w:[ 0 ] /st:0
  or g10 (.I0(A), .I1(B), .Z(w9));   //: @(458,207) /sn:0 /w:[ 7 7 1 ]
  concat g25 (.I0(w3), .I1(w4), .I2(w4), .I3(w4), .I4(w4), .I5(w4), .I6(w4), .I7(w4), .I8(w4), .I9(w4), .I10(w4), .I11(w4), .I12(w4), .I13(w4), .I14(w4), .I15(w4), .I16(w4), .I17(w4), .I18(w4), .I19(w4), .I20(w4), .I21(w4), .I22(w4), .I23(w4), .I24(w4), .I25(w4), .I26(w4), .I27(w4), .I28(w4), .I29(w4), .I30(w4), .I31(w4), .Z(w18));   //: @(778,415) /sn:0 /R:1 /w:[ 1 61 63 65 67 69 71 73 75 77 79 81 83 85 87 89 91 93 95 97 99 101 103 105 107 109 111 113 115 117 119 121 1 ] /dr:0
  //: joint g49 (w4) @(803, 451) /w:[ 38 84 37 -1 ]
  //: joint g6 (A) @(316, 178) /w:[ 2 1 -1 4 ]
  //: joint g50 (w4) @(783, 451) /w:[ 34 88 33 -1 ]
  mux g9 (.I0(w7), .I1(w9), .I2(w2), .I3(!w7), .I4(w13), .I5(w13), .I6(w17), .I7(w18), .S(w0), .Z(ALU_RES));   //: @(703,314) /sn:0 /R:1 /w:[ 3 0 1 5 3 5 3 0 1 0 ] /ss:1 /do:0
  //: joint g7 (B) @(358, 183) /w:[ 2 1 -1 4 ]
  //: joint g35 (w4) @(713, 451) /w:[ 20 102 19 -1 ]
  //: joint g56 (w4) @(663, 451) /w:[ 10 112 9 -1 ]
  //: joint g58 (w4) @(633, 451) /w:[ 4 118 3 -1 ]
  //: joint g22 (w7) @(664, 290) /w:[ 2 1 -1 4 ]
  //: joint g33 (w4) @(673, 451) /w:[ 12 110 11 -1 ]
  //: joint g36 (w4) @(733, 451) /w:[ 24 98 23 -1 ]
  //: joint g41 (w4) @(833, 451) /w:[ 44 78 43 -1 ]
  //: joint g45 (w4) @(893, 451) /w:[ 56 66 55 -1 ]
  //: joint g54 (w4) @(703, 451) /w:[ 18 104 17 -1 ]
  //: joint g40 (w4) @(813, 451) /w:[ 40 82 39 -1 ]
  //: joint g42 (w4) @(853, 451) /w:[ 48 74 47 -1 ]
  //: joint g52 (w4) @(743, 451) /w:[ 26 96 25 -1 ]
  //: joint g12 (B) @(358, 209) /w:[ 6 5 -1 8 ]
  //: joint g34 (w4) @(693, 451) /w:[ 16 106 15 -1 ]
  //: joint g46 (w4) @(863, 451) /w:[ 50 72 49 -1 ]
  //: joint g57 (w4) @(643, 451) /w:[ 6 116 5 -1 ]
  add g5 (.A(B), .B(A), .S(w2), .CI(w5), .CO(w6));   //: @(461,266) /sn:0 /R:1 /w:[ 11 11 0 0 1 ]
  //: joint g11 (A) @(316, 204) /w:[ 6 5 -1 8 ]
  //: joint g14 (A) @(316, 250) /w:[ 10 9 -1 12 ]
  //: joint g19 (w4) @(623, 451) /w:[ 2 120 1 -1 ]
  //: comment g61 /dolink:0 /link:"" @(554,334) /sn:0 /R:2
  //: /line:"unused pins"
  //: /line:"   0011"
  //: /line:"   0100"
  //: /line:"   0101"
  //: /end
  //: joint g21 (w13) @(635, 317) /w:[ 2 -1 1 4 ]
  //: supply0 g20 (w4) @(593,451) /sn:0 /R:3 /w:[ 0 ]
  //: joint g32 (w4) @(653, 451) /w:[ 8 114 7 -1 ]
  //: joint g15 (B) @(358, 282) /w:[ 10 9 -1 12 ]
  //: input g0 (A) @(316,126) /sn:0 /R:3 /w:[ 0 ]
  //: joint g38 (w4) @(773, 451) /w:[ 32 90 31 -1 ]
  //: joint g43 (w4) @(873, 451) /w:[ 52 70 51 -1 ]
  tran g27(.Z(w3), .I(w17[31]));   //: @(564,396) /sn:0 /R:1 /w:[ 0 1 2 ] /ss:1
  //: joint g48 (w4) @(823, 451) /w:[ 42 80 41 -1 ]
  //: joint g37 (w4) @(753, 451) /w:[ 28 94 27 -1 ]
  tran g62(.Z(w0), .I(ALU_OP[2:0]));   //: @(703,248) /sn:0 /R:1 /w:[ 0 2 1 ] /ss:1
  //: joint g55 (w4) @(683, 451) /w:[ 14 108 13 -1 ]
  //: supply0 g13 (w5) @(482,244) /sn:0 /w:[ 1 ]
  //: joint g53 (w4) @(723, 451) /w:[ 22 100 21 -1 ]

endmodule

module BRegs32x32(Read2, Write, Read1, Data2, Data1, clr, clk, RegWrite, WriteData);
//: interface  /sz:(147, 182) /bd:[ Ti0>clr(66/147) Ti1>clr(66/147) Ti2>clr(66/147) Ti3>clr(66/147) Li0>Read1[4:0](32/182) Li1>Read2[4:0](72/182) Li2>Write[4:0](108/182) Li3>WriteData[31:0](148/182) Li4>Read1[4:0](32/182) Li5>Read2[4:0](72/182) Li6>Write[4:0](108/182) Li7>WriteData[31:0](148/182) Li8>WriteData[31:0](148/182) Li9>Write[4:0](108/182) Li10>Read2[4:0](72/182) Li11>Read1[4:0](32/182) Li12>WriteData[31:0](148/182) Li13>Write[4:0](108/182) Li14>Read2[4:0](72/182) Li15>Read1[4:0](32/182) Bi0>clk(108/147) Bi1>RegWrite(40/147) Bi2>clk(108/147) Bi3>RegWrite(40/147) Bi4>RegWrite(40/147) Bi5>clk(108/147) Bi6>RegWrite(40/147) Bi7>clk(108/147) Ro0<Data1[31:0](47/182) Ro1<Data2[31:0](139/182) Ro2<Data1[31:0](47/182) Ro3<Data2[31:0](139/182) Ro4<Data2[31:0](139/182) Ro5<Data1[31:0](47/182) Ro6<Data2[31:0](139/182) Ro7<Data1[31:0](47/182) ]
output [31:0] Data2;    //: /sn:0 {0}(668,485)(668,474)(669,474)(669,464){1}
//: {2}(671,462)(779,462){3}
//: {4}(669,460)(669,445){5}
input [4:0] Write;    //: /sn:0 {0}(-238,-38)(-138,-38)(-138,-37)(-66,-37){1}
//: {2}(-65,-37)(-28,-37){3}
//: {4}(-27,-37)(-16,-37){5}
input [31:0] WriteData;    //: /sn:0 {0}(669,157)(669,124){1}
//: {2}(671,122)(817,122)(817,94){3}
//: {4}(669,120)(669,75)(481,75){5}
//: {6}(477,75)(292,75){7}
//: {8}(288,75)(89,75){9}
//: {10}(85,75)(-104,75)(-104,73)(-237,73){11}
//: {12}(87,77)(87,157){13}
//: {14}(290,77)(290,107)(291,107)(291,152){15}
//: {16}(479,77)(479,157){17}
output [31:0] Data1;    //: /sn:0 {0}(59,382)(59,441){1}
//: {2}(61,443)(204,443)(204,487){3}
//: {4}(59,445)(59,465){5}
supply1 w21;    //: /sn:0 {0}(82,3)(57,3)(57,-11){1}
input clr;    //: /sn:0 {0}(721,193)(731,193)(731,-83)(543,-83){1}
//: {2}(539,-83)(355,-83){3}
//: {4}(351,-83)(150,-83){5}
//: {6}(146,-83)(-44,-83)(-44,-92)(-235,-92){7}
//: {8}(148,-81)(148,193)(139,193){9}
//: {10}(353,-81)(353,188)(343,188){11}
//: {12}(541,-81)(541,193)(531,193){13}
input RegWrite;    //: /sn:0 {0}(-237,263)(-71,263){1}
//: {2}(-67,263)(171,263){3}
//: {4}(175,263)(370,263){5}
//: {6}(374,263)(552,263)(552,219)(556,219){7}
//: {8}(372,261)(372,219)(383,219){9}
//: {10}(173,261)(173,214)(183,214){11}
//: {12}(-69,261)(-69,219)(-38,219){13}
input clk;    //: /sn:0 {0}(556,214)(542,214)(542,285)(364,285){1}
//: {2}(362,283)(362,214)(383,214){3}
//: {4}(360,285)(167,285){5}
//: {6}(165,283)(165,209)(183,209){7}
//: {8}(163,285)(-56,285){9}
//: {10}(-58,283)(-58,214)(-38,214){11}
//: {12}(-60,285)(-237,285){13}
input [4:0] Read1;    //: {0}(-237,96)(-208,96)(-208,95)(-124,95){1}
//: {2}(-123,95)(-96,95){3}
//: {4}(-95,95)(-78,95){5}
input [4:0] Read2;    //: {0}(-237,145)(-141,145){1}
//: {2}(-140,145)(-123,145)(-123,144)(-94,144){3}
//: {4}(-93,144)(-79,144){5}
wire [1:0] w6;    //: /sn:0 {0}(36,369)(-123,369)(-123,99){1}
wire w16;    //: /sn:0 {0}(39,205)(-50,205)(-50,39)(88,39)(88,19){1}
wire w4;    //: /sn:0 {0}(112,19)(112,46)(370,46)(370,205)(431,205){1}
wire [31:0] w3;    //: /sn:0 {0}(77,353)(77,334)(659,334)(659,228){1}
wire [31:0] R2;    //: {0}(65,353)(65,319)(469,319)(469,228){1}
wire [31:0] w0;    //: /sn:0 {0}(651,416)(651,398)(105,398)(105,228){1}
wire w22;    //: /sn:0 {0}(404,217)(431,217){1}
wire w20;    //: /sn:0 {0}(124,19)(124,29)(556,29)(556,205)(621,205){1}
wire [2:0] w19;    //: /sn:0 {0}(431,169)(419,169)(419,109){1}
//: {2}(421,107)(606,107)(606,169)(621,169){3}
//: {4}(417,107)(297,107)(297,106)(231,106){5}
//: {6}(227,106)(25,106){7}
//: {8}(21,106)(-95,106)(-95,99){9}
//: {10}(23,108)(23,169)(39,169){11}
//: {12}(229,108)(229,164)(243,164){13}
wire [2:0] w18;    //: /sn:0 {0}(431,180)(402,180)(402,125){1}
//: {2}(404,123)(589,123)(589,180)(621,180){3}
//: {4}(400,123)(279,123)(279,122)(212,122){5}
//: {6}(208,122)(8,122){7}
//: {8}(4,122)(-93,122)(-93,139){9}
//: {10}(6,124)(6,180)(39,180){11}
//: {12}(210,124)(210,175)(243,175){13}
wire w23;    //: /sn:0 {0}(577,217)(621,217){1}
wire [1:0] w10;    //: /sn:0 {0}(-140,149)(-140,432)(646,432){1}
wire [2:0] w24;    //: /sn:0 {0}(431,193)(381,193)(381,141){1}
//: {2}(383,139)(568,139)(568,193)(621,193){3}
//: {4}(379,139)(260,139)(260,138)(195,138){5}
//: {6}(191,138)(-13,138){7}
//: {8}(-17,138)(-65,138)(-65,-33){9}
//: {10}(-15,140)(-15,193)(39,193){11}
//: {12}(193,140)(193,188)(243,188){13}
wire w31;    //: /sn:0 {0}(243,200)(178,200)(178,60)(100,60)(100,19){1}
wire w1;    //: /sn:0 {0}(-17,217)(39,217){1}
wire [31:0] R1;    //: {0}(281,223)(281,308)(53,308)(53,353){1}
wire [31:0] R3;    //: {0}(687,228)(687,416){1}
wire [1:0] w11;    //: /sn:0 {0}(-27,-33)(-27,-23)(106,-23)(106,-10){1}
wire w2;    //: /sn:0 {0}(243,212)(204,212){1}
wire [31:0] R0;    //: {0}(77,228)(77,299)(41,299)(41,353){1}
wire [31:0] w5;    //: /sn:0 {0}(675,416)(675,372)(497,372)(497,228){1}
wire [31:0] w9;    //: /sn:0 {0}(663,416)(663,387)(309,387)(309,223){1}
//: enddecls

  //: joint g8 (w18) @(6, 122) /w:[ 7 -1 8 10 ]
  //: input g4 (Read2) @(-239,145) /sn:0 /w:[ 0 ]
  //: joint g44 (clr) @(353, -83) /w:[ 3 -1 4 10 ]
  //: input g3 (Write) @(-240,-38) /sn:0 /w:[ 0 ]
  //: joint g16 (clk) @(165, 285) /w:[ 5 6 8 -1 ]
  //: joint g47 (clr) @(541, -83) /w:[ 1 -1 2 12 ]
  //: input g17 (Read1) @(-239,96) /sn:0 /w:[ 0 ]
  //: joint g26 (w19) @(229, 106) /w:[ 5 -1 6 12 ]
  //: output g2 (Data2) @(668,482) /sn:0 /R:3 /w:[ 0 ]
  tran g23(.Z(w24), .I(Write[2:0]));   //: @(-65,-39) /sn:0 /R:1 /w:[ 9 1 2 ] /ss:1
  tran g30(.Z(w10), .I(Read2[4:3]));   //: @(-140,143) /sn:0 /R:1 /w:[ 0 1 2 ] /ss:1
  //: output g1 (Data1) @(59,462) /sn:0 /R:3 /w:[ 5 ]
  //: joint g39 (RegWrite) @(372, 263) /w:[ 6 8 5 -1 ]
  Regs8x32 g24 (.DIN(WriteData), .SD(w24), .SA(w19), .SB(w18), .RegWr(w31), .clk(w2), .clr(clr), .AOUT(R1), .BOUT(w9));   //: @(244, 153) /sz:(98, 69) /sn:0 /p:[ Ti0>15 Li0>13 Li1>13 Li2>13 Li3>0 Li4>0 Ri0>11 Bo0<0 Bo1<1 ]
  Regs8x32 g29 (.DIN(WriteData), .SD(w24), .SA(w19), .SB(w18), .RegWr(w4), .clk(w22), .clr(clr), .AOUT(R2), .BOUT(w5));   //: @(432, 158) /sz:(98, 69) /sn:0 /p:[ Ti0>17 Li0>0 Li1>0 Li2>0 Li3>1 Li4>1 Ri0>13 Bo0<1 Bo1<1 ]
  //: comment g51 /dolink:0 /link:"" @(395,229) /sn:0
  //: /line:"Regs 16-23"
  //: /end
  tran g18(.Z(w19), .I(Read1[2:0]));   //: @(-95,93) /sn:0 /R:1 /w:[ 9 3 4 ] /ss:1
  //: supply1 g10 (w21) @(68,-11) /sn:0 /w:[ 1 ]
  //: joint g25 (w18) @(210, 122) /w:[ 5 -1 6 12 ]
  //: comment g49 /dolink:0 /link:"" @(210,225) /sn:0
  //: /line:"Regs 8-15"
  //: /end
  //: comment g50 /dolink:0 /link:"" @(585,229) /sn:0
  //: /line:"Regs 24-31"
  //: /end
  Regs8x32 g6 (.DIN(WriteData), .SD(w24), .SA(w19), .SB(w18), .RegWr(w16), .clk(w1), .clr(clr), .AOUT(R0), .BOUT(w0));   //: @(40, 158) /sz:(98, 69) /sn:0 /p:[ Ti0>13 Li0>11 Li1>11 Li2>11 Li3>0 Li4>1 Ri0>9 Bo0<0 Bo1<1 ]
  //: joint g7 (w19) @(23, 106) /w:[ 7 -1 8 10 ]
  demux g9 (.I(w11), .E(w21), .Z0(w16), .Z1(w31), .Z2(w4), .Z3(w20));   //: @(106,3) /sn:0 /w:[ 1 0 1 1 0 0 ]
  and g35 (.I0(clk), .I1(RegWrite), .Z(w22));   //: @(394,217) /sn:0 /delay:" 1" /w:[ 3 9 0 ]
  //: joint g56 (Data1) @(59, 443) /w:[ 2 1 -1 4 ]
  tran g31(.Z(w6), .I(Read1[4:3]));   //: @(-123,93) /sn:0 /R:1 /w:[ 1 1 2 ] /ss:1
  tran g22(.Z(w18), .I(Read2[2:0]));   //: @(-93,142) /sn:0 /R:1 /w:[ 9 3 4 ] /ss:0
  and g36 (.I0(clk), .I1(RegWrite), .Z(w23));   //: @(567,217) /sn:0 /delay:" 1" /w:[ 0 7 0 ]
  //: joint g41 (w19) @(419, 107) /w:[ 2 -1 4 1 ]
  //: joint g45 (WriteData) @(479, 75) /w:[ 5 -1 6 16 ]
  and g33 (.I0(clk), .I1(RegWrite), .Z(w1));   //: @(-27,217) /sn:0 /delay:" 1" /w:[ 11 13 0 ]
  led g54 (.I(Data1));   //: @(204,494) /sn:0 /R:2 /w:[ 3 ] /type:2
  //: input g42 (clr) @(-237,-92) /sn:0 /w:[ 7 ]
  //: joint g40 (w18) @(402, 123) /w:[ 2 -1 4 1 ]
  led g52 (.I(WriteData));   //: @(817,87) /sn:0 /w:[ 3 ] /type:2
  //: input g12 (clk) @(-239,285) /sn:0 /w:[ 13 ]
  and g34 (.I0(clk), .I1(RegWrite), .Z(w2));   //: @(194,212) /sn:0 /delay:" 1" /w:[ 7 11 1 ]
  //: joint g28 (w24) @(381, 139) /w:[ 2 -1 4 1 ]
  Regs8x32 g46 (.DIN(WriteData), .SD(w24), .SA(w19), .SB(w18), .RegWr(w20), .clk(w23), .clr(clr), .AOUT(w3), .BOUT(R3));   //: @(622, 158) /sz:(98, 69) /sn:0 /p:[ Ti0>0 Li0>3 Li1>3 Li2>3 Li3>1 Li4>1 Ri0>0 Bo0<1 Bo1<0 ]
  //: joint g57 (Data2) @(669, 462) /w:[ 2 4 -1 1 ]
  //: joint g11 (w24) @(-15, 138) /w:[ 7 -1 8 10 ]
  mux g14 (.I0(R0), .I1(R1), .I2(R2), .I3(w3), .S(w6), .Z(Data1));   //: @(59,369) /sn:0 /w:[ 1 1 0 0 0 0 ] /ss:0 /do:0
  tran g5(.Z(w11), .I(Write[4:3]));   //: @(-27,-39) /sn:0 /R:1 /w:[ 0 3 4 ] /ss:1
  //: joint g19 (clk) @(-58, 285) /w:[ 9 10 12 -1 ]
  //: joint g21 (w24) @(193, 138) /w:[ 5 -1 6 12 ]
  //: input g32 (RegWrite) @(-239,263) /sn:0 /w:[ 0 ]
  //: joint g20 (WriteData) @(87, 75) /w:[ 9 -1 10 12 ]
  //: joint g38 (RegWrite) @(173, 263) /w:[ 4 10 3 -1 ]
  //: joint g15 (clk) @(362, 285) /w:[ 1 2 4 -1 ]
  //: joint g43 (clr) @(148, -83) /w:[ 5 -1 6 8 ]
  //: input g0 (WriteData) @(-239,73) /sn:0 /w:[ 11 ]
  //: joint g27 (WriteData) @(290, 75) /w:[ 7 -1 8 14 ]
  //: comment g48 /dolink:0 /link:"" @(11,228) /sn:0
  //: /line:"Regs 0-7"
  //: /end
  //: joint g37 (RegWrite) @(-69, 263) /w:[ 2 12 1 -1 ]
  //: joint g55 (WriteData) @(669, 122) /w:[ 2 4 -1 1 ]
  mux g13 (.I0(w0), .I1(w9), .I2(w5), .I3(R3), .S(w10), .Z(Data2));   //: @(669,432) /sn:0 /w:[ 0 0 0 1 1 5 ] /ss:0 /do:0
  led g53 (.I(Data2));   //: @(786,462) /sn:0 /R:3 /w:[ 3 ] /type:2

endmodule

module Regs8x32(SB, SA, BOUT, AOUT, clk, clr, RegWr, SD, DIN);
//: interface  /sz:(98, 69) /bd:[ Ti0>DIN[31:0](47/98) Ti1>DIN[31:0](47/98) Ti2>DIN[31:0](47/98) Ti3>DIN[31:0](47/98) Li0>clk(59/69) Li1>RegWr(47/69) Li2>SB[2:0](22/69) Li3>SA[2:0](11/69) Li4>SD[2:0](35/69) Li5>clk(59/69) Li6>RegWr(47/69) Li7>SB[2:0](22/69) Li8>SA[2:0](11/69) Li9>SD[2:0](35/69) Li10>SD[2:0](35/69) Li11>SA[2:0](11/69) Li12>SB[2:0](22/69) Li13>RegWr(47/69) Li14>clk(59/69) Li15>SD[2:0](35/69) Li16>SA[2:0](11/69) Li17>SB[2:0](22/69) Li18>RegWr(47/69) Li19>clk(59/69) Ri0>clr(35/69) Ri1>clr(35/69) Ri2>clr(35/69) Ri3>clr(35/69) Bo0<BOUT[31:0](65/98) Bo1<AOUT[31:0](37/98) Bo2<BOUT[31:0](65/98) Bo3<AOUT[31:0](37/98) Bo4<AOUT[31:0](37/98) Bo5<BOUT[31:0](65/98) Bo6<AOUT[31:0](37/98) Bo7<BOUT[31:0](65/98) ]
input [31:0] DIN;    //: /sn:0 {0}(531,269)(531,318){1}
//: {2}(533,320)(627,320){3}
//: {4}(631,320)(715,320){5}
//: {6}(719,320)(807,320)(807,429){7}
//: {8}(717,322)(717,352){9}
//: {10}(629,322)(629,433){11}
//: {12}(529,320)(435,320){13}
//: {14}(431,320)(342,320){15}
//: {16}(338,320)(264,320){17}
//: {18}(260,320)(181,320)(181,352){19}
//: {20}(262,322)(262,439){21}
//: {22}(340,322)(340,351){23}
//: {24}(433,322)(433,436){25}
//: {26}(531,322)(531,348){27}
output [31:0] BOUT;    //: /sn:0 {0}(516,697)(516,672){1}
input [2:0] SD;    //: /sn:0 {0}(782,138)(852,138)(852,156){1}
supply1 w21;    //: /sn:0 {0}(828,169)(801,169)(801,153){1}
input [2:0] SB;    //: /sn:0 {0}(466,659)(493,659){1}
input RegWr;    //: /sn:0 {0}(48,363)(68,363)(68,378)(82,378){1}
input [2:0] SA;    //: /sn:0 {0}(256,657)(231,657){1}
input clr;    //: /sn:0 /dp:1 {0}(959,337)(1032,337){1}
input clk;    //: /sn:0 {0}(82,383)(68,383)(68,398)(55,398){1}
output [31:0] AOUT;    //: /sn:0 {0}(279,670)(279,702){1}
wire [31:0] w16;    //: /sn:0 {0}(531,369)(531,574)(520,574){1}
//: {2}(516,574)(282,574)(282,641){3}
//: {4}(518,576)(518,587)(519,587)(519,643){5}
wire w7;    //: /sn:0 {0}(472,451)(513,451)(513,405)(848,405)(848,185){1}
wire [31:0] R5;    //: {0}(288,641)(288,586)(525,586){1}
//: {2}(529,586)(629,586)(629,454){3}
//: {4}(527,588)(527,617)(525,617)(525,643){5}
wire w4;    //: /sn:0 {0}(943,337)(906,337){1}
//: {2}(902,337)(767,337){3}
//: {4}(763,337)(588,337){5}
//: {6}(584,337)(390,337){7}
//: {8}(386,337)(231,337)(231,357)(220,357){9}
//: {10}(388,339)(388,356)(379,356){11}
//: {12}(586,339)(586,353)(570,353){13}
//: {14}(765,339)(765,357)(756,357){15}
//: {16}(904,339)(904,417)(865,417){17}
//: {18}(861,417)(675,417){19}
//: {20}(671,417)(489,417){21}
//: {22}(485,417)(302,417)(302,444)(301,444){23}
//: {24}(487,419)(487,441)(472,441){25}
//: {26}(673,419)(673,438)(668,438){27}
//: {28}(863,419)(863,434)(846,434){29}
wire [31:0] R2;    //: {0}(262,641)(262,537){1}
//: {2}(264,535)(499,535)(499,643){3}
//: {4}(262,533)(262,460){5}
wire w0;    //: /sn:0 {0}(770,439)(764,439)(764,481)(579,481){1}
//: {2}(577,479)(577,443)(592,443){3}
//: {4}(575,481)(390,481){5}
//: {6}(388,479)(388,446)(396,446){7}
//: {8}(386,481)(214,481){9}
//: {10}(212,479)(212,449)(225,449){11}
//: {12}(210,481)(125,481)(125,383){13}
//: {14}(127,381)(291,381){15}
//: {16}(295,381)(477,381){17}
//: {18}(481,381)(660,381)(660,362)(680,362){19}
//: {20}(479,379)(479,358)(494,358){21}
//: {22}(293,379)(293,361)(303,361){23}
//: {24}(125,379)(125,362)(144,362){25}
//: {26}(123,381)(103,381){27}
wire w3;    //: /sn:0 {0}(835,185)(835,397)(330,397)(330,454)(301,454){1}
wire [31:0] R7;    //: {0}(807,450)(807,609)(541,609){1}
//: {2}(537,609)(302,609)(302,641){3}
//: {4}(539,611)(539,643){5}
wire w12;    //: /sn:0 {0}(756,367)(787,367)(787,258)(868,258)(868,185){1}
wire w10;    //: /sn:0 {0}(846,444)(875,444)(875,185){1}
wire [31:0] R4;    //: {0}(340,372)(340,545){1}
//: {2}(342,547)(505,547)(505,643){3}
//: {4}(338,547)(268,547)(268,641){5}
wire [31:0] R3;    //: {0}(512,643)(512,559)(435,559){1}
//: {2}(433,557)(433,457){3}
//: {4}(431,559)(275,559)(275,641){5}
wire w8;    //: /sn:0 {0}(220,367)(249,367)(249,213)(828,213)(828,185){1}
wire Z5;    //: /sn:0 {0}(861,185)(861,413)(700,413)(700,448)(668,448){1}
wire w14;    //: /sn:0 {0}(379,366)(414,366)(414,229)(841,229)(841,185){1}
wire [31:0] R0;    //: {0}(492,643)(492,523)(257,523){1}
//: {2}(253,523)(181,523)(181,373){3}
//: {4}(255,525)(255,641){5}
wire w15;    //: /sn:0 {0}(570,363)(608,363)(608,244)(855,244)(855,185){1}
wire [31:0] R10;    //: /sn:0 {0}(295,641)(295,600)(530,600){1}
//: {2}(534,600)(717,600)(717,373){3}
//: {4}(532,602)(532,643){5}
//: enddecls

  //: joint g8 (w16) @(518, 574) /w:[ 1 -1 2 4 ]
  //: input g4 (SB) @(464,659) /sn:0 /w:[ 0 ]
  //: input g3 (SA) @(229,657) /sn:0 /w:[ 1 ]
  //: joint g16 (R3) @(433, 559) /w:[ 1 2 4 -1 ]
  //: joint g17 (R4) @(340, 547) /w:[ 2 1 4 -1 ]
  //: joint g26 (DIN) @(340, 320) /w:[ 15 -1 16 22 ]
  register R5 (.Q(R5), .D(DIN), .EN(Z5), .CLR(w4), .CK(!w0));   //: @(629,443) /w:[ 3 11 1 27 3 ]
  //: output g2 (BOUT) @(516,694) /sn:0 /R:3 /w:[ 0 ]
  //: joint g23 (w4) @(765, 337) /w:[ 3 -1 4 14 ]
  //: joint g30 (w0) @(212, 481) /w:[ 9 10 12 -1 ]
  //: output g1 (AOUT) @(279,699) /sn:0 /R:3 /w:[ 1 ]
  //: joint g39 (DIN) @(262, 320) /w:[ 17 -1 18 20 ]
  //: joint g24 (DIN) @(531, 320) /w:[ 2 1 12 26 ]
  //: joint g29 (w0) @(388, 481) /w:[ 5 6 8 -1 ]
  register R2 (.Q(R4), .D(DIN), .EN(w14), .CLR(w4), .CK(!w0));   //: @(340,361) /w:[ 0 23 0 11 23 ]
  register R7 (.Q(R7), .D(DIN), .EN(w10), .CLR(w4), .CK(!w0));   //: @(807,439) /w:[ 0 7 0 29 0 ]
  //: joint g18 (R2) @(262, 535) /w:[ 2 4 -1 1 ]
  //: supply1 g10 (w21) @(812,153) /sn:0 /w:[ 1 ]
  not g25 (.I(clr), .Z(w4));   //: @(953,337) /sn:0 /R:2 /w:[ 0 0 ]
  //: joint g6 (R7) @(539, 609) /w:[ 1 -1 2 4 ]
  register R6 (.Q(R10), .D(DIN), .EN(w12), .CLR(w4), .CK(!w0));   //: @(717,362) /w:[ 3 9 0 15 19 ]
  //: joint g7 (R10) @(532, 600) /w:[ 2 -1 1 4 ]
  register R4 (.Q(w16), .D(DIN), .EN(w15), .CLR(w4), .CK(!w0));   //: @(531,358) /w:[ 0 27 0 13 21 ]
  demux g9 (.I(SD), .E(w21), .Z0(!w8), .Z1(!w3), .Z2(!w14), .Z3(!w7), .Z4(!w15), .Z5(!Z5), .Z6(!w12), .Z7(!w10));   //: @(852,169) /sn:0 /w:[ 1 0 1 0 1 1 1 0 1 1 ]
  and g35 (.I0(RegWr), .I1(clk), .Z(w0));   //: @(93,381) /sn:0 /delay:" 1" /w:[ 1 0 27 ]
  //: joint g31 (w4) @(863, 417) /w:[ 17 -1 18 28 ]
  //: joint g22 (w4) @(586, 337) /w:[ 5 -1 6 12 ]
  register R3 (.Q(R3), .D(DIN), .EN(w7), .CLR(w4), .CK(!w0));   //: @(433,446) /w:[ 3 25 0 25 7 ]
  register R1 (.Q(R2), .D(DIN), .EN(w3), .CLR(w4), .CK(!w0));   //: @(262,449) /w:[ 5 21 1 23 11 ]
  //: joint g36 (w4) @(904, 337) /w:[ 1 -1 2 16 ]
  //: joint g41 (DIN) @(717, 320) /w:[ 6 -1 5 8 ]
  //: joint g33 (w4) @(673, 417) /w:[ 19 -1 20 26 ]
  //: joint g42 (DIN) @(629, 320) /w:[ 4 -1 3 10 ]
  //: joint g40 (DIN) @(433, 320) /w:[ 13 -1 14 24 ]
  //: joint g12 (w0) @(479, 381) /w:[ 18 20 17 -1 ]
  //: input g34 (clk) @(53,398) /sn:0 /w:[ 1 ]
  //: input g28 (clr) @(1034,337) /sn:0 /R:2 /w:[ 1 ]
  //: joint g11 (w0) @(293, 381) /w:[ 16 22 15 -1 ]
  //: input g5 (RegWr) @(46,363) /sn:0 /w:[ 0 ]
  mux g14 (.I0(R0), .I1(R2), .I2(R4), .I3(R3), .I4(w16), .I5(R5), .I6(R10), .I7(R7), .S(SA), .Z(AOUT));   //: @(279,657) /sn:0 /w:[ 5 0 5 5 3 0 0 3 0 0 ] /ss:0 /do:0
  //: joint g19 (R0) @(255, 523) /w:[ 1 -1 2 4 ]
  //: joint g21 (w4) @(388, 337) /w:[ 7 -1 8 10 ]
  //: joint g32 (w4) @(487, 417) /w:[ 21 -1 22 24 ]
  //: input g20 (SD) @(780,138) /sn:0 /w:[ 0 ]
  register R0 (.Q(R0), .D(DIN), .EN(w8), .CLR(w4), .CK(!w0));   //: @(181,362) /w:[ 3 19 0 9 25 ]
  //: joint g38 (w0) @(577, 481) /w:[ 1 2 4 -1 ]
  //: joint g15 (R5) @(527, 586) /w:[ 2 -1 1 4 ]
  //: input g0 (DIN) @(531,267) /sn:0 /R:3 /w:[ 0 ]
  //: joint g27 (w0) @(125, 381) /w:[ 14 24 26 13 ]
  mux g13 (.I0(R0), .I1(R2), .I2(R4), .I3(R3), .I4(w16), .I5(R5), .I6(R10), .I7(R7), .S(SB), .Z(BOUT));   //: @(516,659) /sn:0 /w:[ 0 3 3 0 5 5 5 5 1 1 ] /ss:0 /do:0

endmodule

module FETCH(clk, PCNew, Reset, Inst, PCNext);
//: interface  /sz:(113, 114) /bd:[ Li0>Reset(33/114) Li1>PCNew[31:0](66/114) Li2>clk(96/114) Li3>Reset(33/114) Li4>PCNew[31:0](66/114) Li5>clk(96/114) Ro0<PCNext[31:0](36/114) Ro1<Inst[31:0](88/114) Ro2<PCNext[31:0](36/114) Ro3<Inst[31:0](88/114) ]
supply0 w6;    //: /sn:0 {0}(521,437)(521,414){1}
supply0 w0;    //: /sn:0 {0}(469,353)(469,326)(454,326)(454,351){1}
input [31:0] PCNew;    //: /sn:0 {0}(383,389)(438,389){1}
output [31:0] Inst;    //: /sn:0 /dp:1 {0}(594,387)(538,387){1}
output [31:0] PCNext;    //: /sn:0 /dp:1 {0}(604,336)(493,336)(493,387){1}
//: {2}(495,389)(503,389){3}
//: {4}(491,389)(459,389){5}
input Reset;    //: /sn:0 {0}(381,328)(444,328)(444,351){1}
input clk;    //: /sn:0 {0}(381,447)(449,447)(449,427){1}
//: enddecls

  //: supply0 g4 (w0) @(469,359) /sn:0 /w:[ 0 ]
  //: input g3 (clk) @(379,447) /sn:0 /w:[ 0 ]
  //: input g2 (PCNew) @(381,389) /sn:0 /w:[ 0 ]
  rom fetch_rom (.A(PCNext), .D(Inst), .OE(w6));   //: @(521,388) /sn:0 /w:[ 3 1 1 ] /mem:"/media/sf_URV/EC/Practica2_EstructuraComputadors/FILES/mult.mem"
  //: input g1 (Reset) @(379,328) /sn:0 /w:[ 0 ]
  //: output g12 (Inst) @(591,387) /sn:0 /w:[ 0 ]
  //: supply0 g11 (w6) @(521,443) /sn:0 /w:[ 0 ]
  register g5 (.Q(PCNext), .D(PCNew), .EN(w0), .CLR(!Reset), .CK(!clk));   //: @(449,389) /sn:0 /R:1 /w:[ 5 1 1 1 1 ]
  //: joint g0 (PCNext) @(493, 389) /w:[ 2 1 4 -1 ]
  //: output g13 (PCNext) @(601,336) /sn:0 /w:[ 0 ]

endmodule

module main;    //: root_module
supply1 w7;    //: /sn:0 {0}(1372,270)(1372,289){1}
wire [7:0] w6;    //: /sn:0 {0}(1351,0)(1361,0){1}
wire [31:0] w13;    //: /sn:0 /dp:1 {0}(502,103)(542,103){1}
//: {2}(544,101)(544,-145)(1081,-145){3}
//: {4}(544,105)(544,207)(452,207){5}
wire [31:0] w16;    //: /sn:0 {0}(452,237)(542,237){1}
//: {2}(546,237)(582,237){3}
//: {4}(584,235)(584,189){5}
//: {6}(584,188)(584,15){7}
//: {8}(584,14)(584,-163){9}
//: {10}(584,-164)(584,-175){11}
//: {12}(584,239)(584,263){13}
//: {14}(584,264)(584,287){15}
//: {16}(584,288)(584,378){17}
//: {18}(584,379)(584,392){19}
//: {20}(544,239)(544,335)(526,335){21}
wire [31:0] Data2;    //: /sn:0 /dp:1 {0}(1195,227)(1175,227)(1175,327){1}
//: {2}(1177,329)(1358,329){3}
//: {4}(1175,331)(1175,341)(920,341){5}
//: {6}(916,341)(865,341)(865,293){7}
//: {8}(867,291)(878,291){9}
//: {10}(879,291)(921,291){11}
//: {12}(863,291)(848,291){13}
//: {14}(918,343)(918,450)(928,450){15}
wire w34;    //: /sn:0 {0}(879,76)(902,76){1}
//: {2}(906,76)(916,76){3}
//: {4}(904,78)(904,145)(814,145){5}
wire w39;    //: /sn:0 {0}(1459,107)(804,107)(804,93){1}
wire w25;    //: /sn:0 {0}(1351,17)(1361,17){1}
wire [4:0] w4;    //: /sn:0 /dp:1 {0}(588,264)(669,264){1}
//: {2}(673,264)(718,264){3}
//: {4}(671,262)(671,245){5}
wire [31:0] readData;    //: /sn:0 /dp:1 {0}(1358,297)(1332,297)(1332,188){1}
//: {2}(1334,186)(1386,186){3}
//: {4}(1390,186)(1406,186){5}
//: {6}(1388,184)(1388,147)(1490,147){7}
//: {8}(1330,186)(1297,186){9}
wire [4:0] Write;    //: /sn:0 /dp:1 {0}(718,288)(673,288){1}
//: {2}(669,288)(588,288){3}
//: {4}(671,290)(671,299){5}
wire w36;    //: /sn:0 {0}(1361,33)(1351,33){1}
wire [7:0] w22;    //: /sn:0 {0}(1361,8)(1351,8){1}
wire w0;    //: /sn:0 {0}(337,267)(320,267)(320,316){1}
//: {2}(322,318)(336,318){3}
//: {4}(318,318)(200,318){5}
//: {6}(320,320)(320,438)(765,438)(765,417){7}
wire w3;    //: /sn:0 {0}(879,19)(940,19){1}
//: {2}(944,19)(1247,19)(1247,152){3}
//: {4}(942,17)(942,9)(953,9){5}
wire [31:0] w20;    //: /sn:0 /dp:1 {0}(718,347)(686,347)(686,427)(1447,427)(1447,399){1}
//: {2}(1449,397)(1509,397){3}
//: {4}(1447,395)(1447,373){5}
wire w30;    //: /sn:0 {0}(879,-96)(942,-96){1}
//: {2}(946,-96)(1049,-96)(1049,-197)(1155,-197)(1155,-190){3}
//: {4}(944,-98)(944,-108)(954,-108){5}
wire w29;    //: /sn:0 {0}(879,-73)(941,-73){1}
//: {2}(945,-73)(1111,-73){3}
//: {4}(943,-75)(943,-86)(954,-86){5}
wire [25:0] Inm26;    //: /sn:0 /dp:1 {0}(588,-163)(716,-163){1}
//: {2}(720,-163)(1081,-163){3}
//: {4}(718,-165)(718,-191)(433,-191)(433,-180){5}
wire w37;    //: /sn:0 {0}(1351,41)(1361,41){1}
wire [15:0] w19;    //: /sn:0 {0}(708,93)(708,119)(564,119)(564,399){1}
//: {2}(566,401)(673,401)(673,381){3}
//: {4}(675,379)(718,379){5}
//: {6}(671,379)(641,379){7}
//: {8}(640,379)(588,379){9}
//: {10}(562,401)(505,401){11}
wire [31:0] w18;    //: /sn:0 {0}(1084,298)(1143,298){1}
//: {2}(1147,298)(1307,298)(1307,225){3}
//: {4}(1309,223)(1490,223){5}
//: {6}(1307,221)(1307,206)(1406,206){7}
//: {8}(1145,296)(1145,184)(1195,184){9}
wire w12;    //: /sn:0 /dp:1 {0}(879,56)(998,56){1}
//: {2}(1002,56)(1120,56)(1120,83){3}
//: {4}(1000,58)(1000,69)(990,69){5}
wire w10;    //: /sn:0 {0}(1132,-70)(1148,-70)(1148,-76){1}
//: {2}(1150,-78)(1165,-78){3}
//: {4}(1148,-80)(1148,-102){5}
wire w23;    //: /sn:0 /dp:1 {0}(1247,255)(1247,264)(1159,264)(1159,-50)(946,-50){1}
//: {2}(944,-52)(944,-60)(954,-60){3}
//: {4}(942,-50)(879,-50){5}
wire [31:0] Data1;    //: /sn:0 {0}(848,253)(952,253){1}
//: {2}(956,253)(983,253){3}
//: {4}(954,255)(954,352)(1010,352)(1010,359){5}
wire [31:0] SignExtOut;    //: /sn:0 {0}(848,376)(893,376)(893,313){1}
//: {2}(895,311)(921,311){3}
//: {4}(893,309)(893,-122)(939,-122){5}
//: {6}(943,-122)(1081,-122){7}
//: {8}(941,-124)(941,-174){9}
wire w24;    //: /sn:0 {0}(811,417)(811,476){1}
//: {2}(813,478)(1283,478)(1283,255){3}
//: {4}(809,478)(275,478)(275,206){5}
//: {6}(277,204)(337,204){7}
//: {8}(275,202)(275,188){9}
//: {10}(273,204)(249,204){11}
wire [31:0] w21;    //: /sn:0 /dp:1 {0}(1387,313)(1435,313){1}
//: {2}(1439,313)(1491,313){3}
//: {4}(1437,315)(1437,344){5}
wire [5:0] w1;    //: /sn:0 {0}(641,374)(641,80){1}
//: {2}(641,76)(641,48)(687,48){3}
//: {4}(639,78)(631,78){5}
wire w31;    //: /sn:0 {0}(879,-116)(899,-116)(899,-134){1}
//: {2}(901,-136)(907,-136)(907,-136)(910,-136){3}
//: {4}(899,-138)(899,-173)(566,-173)(566,326)(718,326){5}
wire w32;    //: /sn:0 {0}(1361,25)(1351,25){1}
wire w8;    //: /sn:0 {0}(1031,88)(1031,130){1}
//: {2}(1033,132)(1049,132)(1049,62)(1115,62)(1115,83){3}
//: {4}(1029,132)(879,132)(879,286){5}
wire w27;    //: /sn:0 {0}(879,-26)(941,-26){1}
//: {2}(945,-26)(1422,-26)(1422,173){3}
//: {4}(943,-28)(943,-36)(954,-36){5}
wire w17;    //: /sn:0 {0}(1084,255)(1099,255)(1099,161){1}
//: {2}(1099,157)(1099,-68)(1111,-68){3}
//: {4}(1097,159)(1078,159)(1078,147){5}
wire w28;    //: /sn:0 {0}(1372,337)(1372,347){1}
wire w33;    //: /sn:0 {0}(793,147)(780,147)(780,160){1}
wire w35;    //: /sn:0 {0}(1117,104)(1117,148){1}
//: {2}(1115,150)(814,150){3}
//: {4}(1117,152)(1117,360)(1424,360){5}
wire [31:0] w14;    //: /sn:0 /dp:1 {0}(1457,344)(1457,196)(1435,196){1}
wire [4:0] w11;    //: /sn:0 {0}(588,189)(669,189){1}
//: {2}(673,189)(718,189){3}
//: {4}(671,187)(671,175){5}
wire [5:0] w2;    //: /sn:0 {0}(588,15)(656,15){1}
//: {2}(660,15)(687,15){3}
//: {4}(658,13)(658,-15){5}
wire [31:0] w15;    //: /sn:0 /dp:1 {0}(983,301)(950,301){1}
wire w38;    //: /sn:0 {0}(1357,123)(752,123)(752,93){1}
wire [31:0] w5;    //: /sn:0 /dp:1 {0}(337,237)(315,237)(315,-17){1}
//: {2}(317,-19)(343,-19){3}
//: {4}(315,-21)(315,-231)(1354,-231)(1354,-147)(1187,-147){5}
wire [3:0] w26;    //: /sn:0 /dp:1 {0}(879,-2)(1019,-2)(1019,175){1}
//: {2}(1017,177)(995,177){3}
//: {4}(1019,179)(1019,232){5}
wire w9;    //: /sn:0 {0}(879,35)(937,35)(937,40){1}
//: {2}(939,42)(953,42){3}
//: {4}(937,44)(937,278){5}
//: enddecls

  led g75 (.I(w19));   //: @(498,401) /sn:0 /R:1 /w:[ 11 ] /type:2
  //: joint g44 (w29) @(943, -73) /w:[ 2 4 1 -1 ]
  JUMP g4 (.Jump(w30), .SignExt(SignExtOut), .Inm26(Inm26), .PCNext(w13), .PCSrc(w10), .PCin(w5));   //: @(1082, -189) /sz:(104, 86) /sn:0 /p:[ Ti0>3 Li0>7 Li1>3 Li2>3 Bi0>5 Ro0<5 ]
  //: joint g8 (w2) @(658, 15) /w:[ 2 4 1 -1 ]
  //: joint g16 (Write) @(671, 288) /w:[ 1 -1 2 4 ]
  //: comment g47 /dolink:0 /link:"" @(600,42) /sn:0
  //: /line:"funct"
  //: /end
  FETCH g3 (.Reset(w24), .PCNew(w5), .clk(w0), .PCNext(w13), .Inst(w16));   //: @(338, 171) /sz:(113, 114) /sn:0 /p:[ Li0>7 Li1>0 Li2>0 Ro0<5 Ro1<0 ]
  led g109 (.I(w16));   //: @(519,335) /sn:0 /R:1 /w:[ 21 ] /type:2
  //: comment g90 /dolink:0 /link:"" @(1049,394) /sn:0
  //: /line:"Data 1"
  //: /end
  led g26 (.I(w29));   //: @(961,-86) /sn:0 /R:3 /w:[ 5 ] /type:0
  tran g17(.Z(w19), .I(w16[15:0]));   //: @(582,379) /sn:0 /R:2 /w:[ 9 18 17 ] /ss:1
  //: joint g2 (w24) @(275, 204) /w:[ 6 8 10 5 ]
  //: comment g74 /dolink:0 /link:"" @(662,336) /sn:0
  //: /line:"rd"
  //: /end
  led g30 (.I(w27));   //: @(961,-36) /sn:0 /R:3 /w:[ 5 ] /type:0
  led g23 (.I(w30));   //: @(961,-108) /sn:0 /R:3 /w:[ 5 ] /type:0
  //: joint g91 (w24) @(811, 478) /w:[ 2 1 4 -1 ]
  add g92 (.A(!Data2), .B(readData), .S(w21), .CI(w7), .CO(w28));   //: @(1374,313) /sn:0 /R:1 /w:[ 3 0 0 1 0 ]
  //: joint g39 (w34) @(904, 76) /w:[ 2 -1 1 4 ]
  led g86 (.I(Data2));   //: @(935,450) /sn:0 /R:3 /w:[ 15 ] /type:2
  //: comment g77 /dolink:0 /link:"" @(453,367) /sn:0
  //: /line:"Inm16"
  //: /end
  //: joint g24 (Data2) @(865, 291) /w:[ 8 -1 12 7 ]
  clock g1 (.Z(w0));   //: @(187,318) /sn:0 /w:[ 5 ] /omega:3000 /phi:0 /duty:50
  or g104 (.I0(w35), .I1(w34), .Z(w33));   //: @(803,147) /sn:0 /R:2 /w:[ 3 5 0 ]
  //: comment g111 /dolink:0 /link:"" @(422,301) /sn:0
  //: /line:"Instruction"
  //: /end
  //: joint g110 (w16) @(544, 237) /w:[ 2 -1 1 20 ]
  led g60 (.I(w18));   //: @(1497,223) /sn:0 /R:3 /w:[ 5 ] /type:2
  led g29 (.I(w23));   //: @(961,-60) /sn:0 /R:3 /w:[ 3 ] /type:0
  //: comment g51 /dolink:0 /link:"" @(397,65) /sn:0
  //: /line:"PC actual"
  //: /end
  //: joint g82 (SignExtOut) @(941, -122) /w:[ 6 8 5 -1 ]
  //: joint g70 (w4) @(671, 264) /w:[ 2 4 1 -1 ]
  tran g18(.Z(w11), .I(w16[25:21]));   //: @(582,189) /sn:0 /R:2 /w:[ 0 5 6 ] /ss:1
  //: comment g65 /dolink:0 /link:"" @(1544,108) /sn:0
  //: /line:"READ DATA"
  //: /end
  mux g25 (.I0(Data2), .I1(SignExtOut), .S(w9), .Z(w15));   //: @(937,301) /sn:0 /R:1 /w:[ 11 3 5 1 ] /ss:1 /do:1
  led g10 (.I(w1));   //: @(624,78) /sn:0 /R:1 /w:[ 5 ] /type:2
  mux g94 (.I0(w14), .I1(w21), .S(w35), .Z(w20));   //: @(1447,360) /sn:0 /w:[ 0 5 5 5 ] /ss:0 /do:1
  //: comment g103 /dolink:0 /link:"" @(1510,279) /sn:0
  //: /line:"MEM[$b + label] - $a"
  //: /end
  //: joint g64 (Data2) @(1175, 329) /w:[ 2 1 -1 4 ]
  led MEMb__label__a (.I(w21));   //: @(1498,313) /sn:0 /R:3 /w:[ 3 ] /type:2
  //: joint g107 (w20) @(1447, 397) /w:[ 2 4 -1 1 ]
  //: comment g72 /dolink:0 /link:"" @(667,125) /sn:0
  //: /line:"rs"
  //: /end
  led g49 (.I(w13));   //: @(495,103) /sn:0 /R:1 /w:[ 0 ] /type:2
  //: joint g50 (w13) @(544, 103) /w:[ -1 2 1 4 ]
  led g6 (.I(w2));   //: @(658,-22) /sn:0 /w:[ 5 ] /type:2
  //: comment g73 /dolink:0 /link:"" @(668,196) /sn:0
  //: /line:"rt"
  //: /end
  led g68 (.I(w11));   //: @(671,168) /sn:0 /w:[ 5 ] /type:2
  //: joint g58 (w0) @(320, 318) /w:[ 2 1 4 6 ]
  //: joint g56 (w10) @(1148, -78) /w:[ 2 4 -1 1 ]
  and g7 (.I0(w29), .I1(w17), .Z(w10));   //: @(1122,-70) /sn:0 /w:[ 3 3 0 ]
  MEM g9 (.MemWrite(w3), .WriteData(Data2), .Adress(w18), .clk(w24), .MemRead(w23), .ReadData(readData));   //: @(1196, 153) /sz:(100, 101) /sn:0 /p:[ Ti0>3 Li0>0 Li1>9 Bi0>3 Bi1>0 Ro0<9 ]
  //: switch g35 (w24) @(232,204) /sn:0 /w:[ 11 ] /st:0
  //: joint g71 (w11) @(671, 189) /w:[ 2 4 1 -1 ]
  led g59 (.I(w24));   //: @(275,181) /sn:0 /w:[ 9 ] /type:0
  led g31 (.I(w3));   //: @(960,9) /sn:0 /R:3 /w:[ 5 ] /type:0
  //: joint g22 (w31) @(899, -136) /w:[ 2 4 -1 1 ]
  //: joint g98 (w12) @(1000, 56) /w:[ 2 -1 1 4 ]
  //: joint g102 (w18) @(1307, 223) /w:[ 4 6 -1 3 ]
  //: joint g87 (Data2) @(918, 341) /w:[ 5 -1 6 14 ]
  led g85 (.I(Data1));   //: @(1010,366) /sn:0 /R:2 /w:[ 5 ] /type:2
  led g67 (.I(Write));   //: @(671,306) /sn:0 /R:2 /w:[ 5 ] /type:2
  //: comment g83 /dolink:0 /link:"" @(913,-224) /sn:0
  //: /line:"SignExtend"
  //: /end
  //: supply1 g99 (w7) @(1383,270) /sn:0 /w:[ 0 ]
  //: comment g36 /dolink:0 /link:"" @(965,207) /sn:0
  //: /line:"ALU OP"
  //: /end
  //: joint g54 (w17) @(1099, 159) /w:[ -1 2 4 1 ]
  //: joint g45 (w30) @(944, -96) /w:[ 2 4 1 -1 ]
  //: joint g41 (w3) @(942, 19) /w:[ 2 4 1 -1 ]
  led g33 (.I(w9));   //: @(960,42) /sn:0 /R:3 /w:[ 3 ] /type:0
  led g81 (.I(SignExtOut));   //: @(941,-181) /sn:0 /w:[ 9 ] /type:2
  led g69 (.I(w4));   //: @(671,238) /sn:0 /w:[ 5 ] /type:2
  //: joint g52 (w5) @(315, -19) /w:[ 2 4 -1 1 ]
  //: joint g42 (w27) @(943, -26) /w:[ 2 4 1 -1 ]
  //: joint g40 (w9) @(937, 42) /w:[ 2 1 -1 4 ]
  //: comment g66 /dolink:0 /link:"" @(408,-56) /sn:0
  //: /line:"PC NEXT"
  //: /end
  led g12 (.I(w26));   //: @(988,177) /sn:0 /R:1 /w:[ 3 ] /type:2
  //: comment g108 /dolink:0 /link:"" @(1561,365) /sn:0
  //: /line:"WriteData"
  //: /end
  led g57 (.I(w0));   //: @(343,318) /sn:0 /R:3 /w:[ 3 ] /type:0
  //: comment g46 /dolink:0 /link:"" @(654,-69) /sn:0
  //: /line:"op"
  //: /end
  mux g28 (.I0(w18), .I1(readData), .S(w27), .Z(w14));   //: @(1422,196) /sn:0 /R:1 /w:[ 7 5 3 1 ] /ss:1 /do:0
  tran g34(.Z(w2), .I(w16[31:26]));   //: @(582,15) /sn:0 /R:2 /w:[ 0 7 8 ] /ss:1
  led g106 (.I(w20));   //: @(1516,397) /sn:0 /R:3 /w:[ 3 ] /type:2
  //: joint g84 (w16) @(584, 237) /w:[ -1 4 3 12 ]
  //: joint g11 (w1) @(641, 78) /w:[ -1 2 4 1 ]
  //: joint g14 (w26) @(1019, 177) /w:[ -1 1 2 4 ]
  tran g5(.Z(w1), .I(w19[5:0]));   //: @(641,377) /sn:0 /R:1 /w:[ 0 8 7 ] /ss:0
  //: joint g96 (w8) @(1031, 132) /w:[ 2 1 4 -1 ]
  tran g112(.Z(w8), .I(Data2[31]));   //: @(879,289) /sn:0 /R:1 /w:[ 5 9 10 ] /ss:0
  tty g114 (.TD(w6), .RD(w22), .RTS(w25), .CTS(w32), .DSR(w36), .DTR(w37));   //: @(1314,22) /sn:0 /w:[ 0 1 0 1 1 0 ]
  led g21 (.I(w31));   //: @(917,-136) /sn:0 /R:3 /w:[ 3 ] /type:0
  tran g19(.Z(w4), .I(w16[20:16]));   //: @(582,264) /sn:0 /R:2 /w:[ 0 14 13 ] /ss:1
  //: joint g61 (readData) @(1332, 186) /w:[ 2 -1 8 1 ]
  //: comment g79 /dolink:0 /link:"" @(421,-135) /sn:0
  //: /line:"Inm26"
  //: /end
  led g78 (.I(Inm26));   //: @(433,-173) /sn:0 /R:2 /w:[ 5 ] /type:2
  tran g20(.Z(Write), .I(w16[15:11]));   //: @(582,288) /sn:0 /R:2 /w:[ 3 16 15 ] /ss:1
  //: joint g32 (w18) @(1145, 298) /w:[ 2 8 1 -1 ]
  //: joint g113 (w19) @(564, 401) /w:[ 2 1 10 -1 ]
  led g63 (.I(readData));   //: @(1497,147) /sn:0 /R:3 /w:[ 7 ] /type:2
  //: joint g100 (readData) @(1388, 186) /w:[ 4 6 3 -1 ]
  and g93 (.I0(w12), .I1(w8), .Z(w35));   //: @(1117,94) /sn:0 /R:3 /w:[ 3 3 0 ]
  led g97 (.I(w12));   //: @(983,69) /sn:0 /R:1 /w:[ 5 ] /type:0
  //: joint g105 (w35) @(1117, 150) /w:[ -1 1 2 4 ]
  //: comment g89 /dolink:0 /link:"" @(1099,446) /sn:0
  //: /line:"Data2"
  //: /end
  //: joint g43 (w23) @(944, -50) /w:[ 1 2 4 -1 ]
  CONTROL g38 (.funct(w1), .op(w2), .label(w19), .WriteTTY(w39), .ReadTTY(w38), .nsubm(w12), .MemWrite(w3), .RegDst(w31), .Jump(w30), .Branch(w29), .MemRead(w23), .MemToReg(w27), .ALUOp(w26), .ALUSrc(w9), .RegWrite(w34));   //: @(688, -139) /sz:(190, 231) /sn:0 /p:[ Li0>3 Li1>3 Bi0>0 Bo0<1 Bo1<1 Ro0<0 Ro1<0 Ro2<0 Ro3<0 Ro4<0 Ro5<5 Ro6<0 Ro7<0 Ro8<0 Ro9<0 ]
  READ g0 (.RegWrite(w33), .SignExtIn(w19), .WriteData(w20), .RegDst(w31), .Write(Write), .Read2(w4), .Read1(w11), .clr(w24), .clk(w0), .SignExtOut(SignExtOut), .Data2(Data2), .Data1(Data1));   //: @(719, 161) /sz:(128, 255) /sn:0 /p:[ Ti0>1 Li0>5 Li1>0 Li2>5 Li3>0 Li4>3 Li5>3 Bi0>0 Bi1>7 Ro0<0 Ro1<13 Ro2<0 ]
  tran g15(.Z(Inm26), .I(w16[25:0]));   //: @(582,-163) /sn:0 /R:2 /w:[ 0 9 10 ] /ss:1
  //: joint g101 (w21) @(1437, 313) /w:[ 2 -1 1 4 ]
  led g48 (.I(w5));   //: @(350,-19) /sn:0 /R:3 /w:[ 3 ] /type:2
  //: joint g27 (SignExtOut) @(893, 311) /w:[ 2 4 -1 1 ]
  //: comment g62 /dolink:0 /link:"" @(1551,192) /sn:0
  //: /line:"ALU RESULT"
  //: /end
  led g37 (.I(w34));   //: @(923,76) /sn:0 /R:3 /w:[ 3 ] /type:0
  //: joint g88 (Data1) @(954, 253) /w:[ 2 -1 1 4 ]
  //: joint g80 (Inm26) @(718, -163) /w:[ 2 4 1 -1 ]
  led g55 (.I(w10));   //: @(1172,-78) /sn:0 /R:3 /w:[ 3 ] /type:0
  led g95 (.I(w8));   //: @(1031,81) /sn:0 /w:[ 0 ] /type:0
  //: joint g76 (w19) @(673, 379) /w:[ 4 -1 6 3 ]
  led g53 (.I(w17));   //: @(1078,140) /sn:0 /w:[ 5 ] /type:0
  ALU g13 (.ALU_OP(w26), .B(w15), .A(Data1), .ALU_RES(w18), .Zero(w17));   //: @(984, 233) /sz:(99, 90) /sn:0 /p:[ Ti0>5 Li0>0 Li1>3 Ro0<0 Ro1<0 ]

endmodule
