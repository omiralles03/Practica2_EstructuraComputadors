//: version "1.8.7"

module Zero(o, i);
//: interface  /sz:(40, 40) /bd:[ Li0>i[31:0](21/40) Ro0<o(22/40) ]
input [31:0] i;    //: /sn:0 {0}(441,304)(494,304){1}
output o;    //: /sn:0 /dp:1 {0}(645,292)(645,317)(802,317){1}
wire w0;    //: /sn:0 {0}(632,194)(645,194)(645,244){1}
wire [31:0] w1;    //: /sn:0 /dp:1 {0}(496,228)(496,252)(631,252){1}
wire [31:0] w5;    //: /sn:0 /dp:1 {0}(660,268)(787,268)(787,239){1}
wire [31:0] w9;    //: /sn:0 {0}(568,303)(602,303)(602,284)(631,284){1}
//: enddecls

  led g4 (.I(w5));   //: @(787,232) /sn:0 /w:[ 1 ] /type:3
  //: dip g3 (w1) @(496,218) /sn:0 /w:[ 0 ] /st:0
  //: switch g2 (w0) @(615,194) /sn:0 /w:[ 0 ] /st:0
  //: output g1 (o) @(799,317) /sn:0 /w:[ 1 ]
  Ca2 g6 (.in(i), .out(w9));   //: @(495, 282) /sz:(72, 40) /sn:0 /p:[ Li0>1 Ro0<0 ]
  add g5 (.A(w9), .B(w1), .S(w5), .CI(w0), .CO(o));   //: @(647,268) /sn:0 /R:1 /w:[ 1 1 0 1 0 ]
  //: input g0 (i) @(439,304) /sn:0 /w:[ 0 ]

endmodule

module Ca2(out, in);
//: interface  /sz:(72, 40) /bd:[ Li0>in[31:0](22/40) Ro0<out[31:0](21/40) ]
input [31:0] in;    //: /sn:0 {0}(494,347)(552,347){1}
supply0 w0;    //: /sn:0 {0}(551,307)(551,297)(566,297)(566,339){1}
output [31:0] out;    //: /sn:0 /dp:1 {0}(581,363)(639,363){1}
wire [31:0] w1;    //: /sn:0 /dp:1 {0}(484,393)(484,379)(552,379){1}
wire w2;    //: /sn:0 /dp:1 {0}(581,419)(581,429)(566,429)(566,387){1}
//: enddecls

  //: supply0 g4 (w0) @(551,313) /sn:0 /w:[ 0 ]
  //: dip g3 (w1) @(484,404) /sn:0 /R:2 /w:[ 0 ] /st:1
  add g2 (.A(w1), .B(in), .S(out), .CI(w0), .CO(w2));   //: @(568,363) /sn:0 /R:1 /w:[ 1 1 0 1 1 ]
  //: output g1 (out) @(636,363) /sn:0 /w:[ 1 ]
  led g5 (.I(w2));   //: @(581,412) /sn:0 /w:[ 0 ] /type:0
  //: input g0 (in) @(492,347) /sn:0 /w:[ 0 ]

endmodule

module ALU(Result, Zero, B, A, ALU_OP);
//: interface  /sz:(94, 87) /bd:[ Ti0>ALU_OP[3:0](45/94) Li0>A[31:0](30/87) Li1>B[31:0](70/87) Ro0<Zero(32/87) Ro1<Result[31:0](66/87) ]
input [31:0] B;    //: /sn:0 /dp:1 {0}(571,193)(270,193)(270,280){1}
//: {2}(272,282)(576,282){3}
//: {4}(270,284)(270,358){5}
//: {6}(268,360)(131,360)(131,153){7}
//: {8}(270,362)(270,411){9}
//: {10}(268,413)(222,413){11}
//: {12}(270,415)(270,454){13}
//: {14}(272,456)(569,456){15}
//: {16}(270,458)(270,599)(446,599){17}
output Zero;    //: /sn:0 {0}(1411,566)(1505,566){1}
input [31:0] A;    //: /sn:0 {0}(317,322)(359,322){1}
//: {2}(361,320)(361,279){3}
//: {4}(363,277)(576,277){5}
//: {6}(361,275)(361,188)(571,188){7}
//: {8}(361,324)(361,344){9}
//: {10}(363,346)(513,346)(513,112){11}
//: {12}(361,348)(361,422){13}
//: {14}(363,424)(569,424){15}
//: {16}(361,426)(361,566)(570,566){17}
output [31:0] Result;    //: /sn:0 /dp:1 {0}(1084,348)(1317,348){1}
//: {2}(1321,348)(1415,348){3}
//: {4}(1319,350)(1319,565)(1369,565){5}
input [3:0] ALU_OP;    //: /sn:0 /dp:1 {0}(1071,325)(1071,123)(1007,123){1}
wire w16;    //: /sn:0 {0}(584,606)(584,636)(610,636)(610,626){1}
wire [31:0] w13;    //: /sn:0 {0}(1011,532)(1011,503){1}
//: {2}(1013,501)(1162,501)(1162,493){3}
//: {4}(1011,499)(1011,346)(1055,346){5}
wire [31:0] w6;    //: /sn:0 /dp:1 {0}(1021,699)(1021,561){1}
wire [31:0] w0;    //: /sn:0 {0}(520,598)(570,598){1}
wire w22;    //: /sn:0 {0}(545,525)(584,525)(584,558){1}
wire [31:0] w3;    //: /sn:0 /dp:1 {0}(1055,328)(710,328)(710,440)(658,440){1}
//: {2}(654,440)(598,440){3}
//: {4}(656,442)(656,476)(801,476)(801,536)(855,536)(855,704)(681,704)(681,694){5}
wire [31:0] w20;    //: /sn:0 {0}(953,644)(953,607)(964,607){1}
//: {2}(968,607)(1001,607)(1001,561){3}
//: {4}(966,605)(966,468)(956,468){5}
//: {6}(954,466)(954,374)(1055,374){7}
//: {8}(952,468)(940,468){9}
//: {10}(938,466)(938,370)(1055,370){11}
//: {12}(936,468)(922,468){13}
//: {14}(920,466)(920,367)(1055,367){15}
//: {16}(918,468)(903,468){17}
//: {18}(901,466)(901,363)(1055,363){19}
//: {20}(899,468)(882,468){21}
//: {22}(880,466)(880,360)(1055,360){23}
//: {24}(878,468)(864,468){25}
//: {26}(862,466)(862,356)(1055,356){27}
//: {28}(860,468)(838,468){29}
//: {30}(836,466)(836,353)(1055,353){31}
//: {32}(834,468)(813,468){33}
//: {34}(811,466)(811,349)(1055,349){35}
//: {36}(809,468)(794,468){37}
//: {38}(792,466)(792,339)(1055,339){39}
//: {40}(790,468)(770,468){41}
//: {42}(768,466)(768,335)(1055,335){43}
//: {44}(766,468)(732,468)(732,332)(1055,332){45}
wire w23;    //: /sn:0 {0}(537,372)(583,372)(583,416){1}
wire w21;    //: /sn:0 {0}(583,464)(583,498)(600,498)(600,488){1}
wire [31:0] w1;    //: /sn:0 /dp:1 {0}(1055,321)(716,321)(716,191)(592,191){1}
wire [31:0] w2;    //: /sn:0 /dp:1 {0}(1055,325)(689,325)(689,280)(597,280){1}
wire w11;    //: /sn:0 {0}(697,545)(988,545){1}
wire [31:0] w9;    //: /sn:0 /dp:3 {0}(599,582)(693,582)(693,545){1}
//: {2}(693,544)(693,342)(1055,342){3}
//: enddecls

  led g44 (.I(A));   //: @(513,105) /sn:0 /w:[ 11 ] /type:3
  //: output g4 (Result) @(1412,348) /sn:0 /w:[ 3 ]
  add g8 (.A(w0), .B(A), .S(w9), .CI(w22), .CO(w16));   //: @(586,582) /sn:0 /R:1 /w:[ 1 17 0 1 0 ]
  //: joint g47 (w3) @(656, 440) /w:[ 1 -1 2 4 ]
  //: output g3 (Zero) @(1502,566) /sn:0 /w:[ 1 ]
  //: joint g16 (B) @(270, 282) /w:[ 2 1 -1 4 ]
  //: joint g17 (B) @(270, 413) /w:[ -1 9 10 12 ]
  led g26 (.I(w13));   //: @(1162,486) /sn:0 /w:[ 3 ] /type:3
  //: input g2 (B) @(220,413) /sn:0 /w:[ 11 ]
  //: comment g23 /dolink:0 /link:"" @(1052,527) /sn:0
  //: /line:"if (A < B)   // bit 31 = 1"
  //: /line:"   ALU = 1;"
  //: /line:"else         // bit 31 = 0"
  //: /line:"   ALU = 0;"
  //: /end
  //: joint g30 (Result) @(1319, 348) /w:[ 2 -1 1 4 ]
  //: input g1 (A) @(315,322) /sn:0 /w:[ 0 ]
  //: dip g24 (w6) @(1021,710) /sn:0 /R:2 /w:[ 0 ] /st:1
  //: joint g39 (w20) @(811, 468) /w:[ 33 34 36 -1 ]
  Zero g29 (.i(Result), .o(Zero));   //: @(1370, 544) /sz:(40, 40) /sn:0 /p:[ Li0>5 Ro0<0 ]
  //: joint g18 (B) @(270, 456) /w:[ 14 13 -1 16 ]
  //: switch g10 (w22) @(528,525) /sn:0 /w:[ 0 ] /st:0
  //: dip g25 (w20) @(953,655) /sn:0 /R:2 /w:[ 0 ] /st:0
  or g6 (.I0(A), .I1(B), .Z(w2));   //: @(587,280) /sn:0 /w:[ 5 3 1 ]
  add g9 (.A(B), .B(A), .S(w3), .CI(w23), .CO(w21));   //: @(585,440) /sn:0 /R:1 /w:[ 15 15 3 1 0 ]
  mux g7 (.I0(w1), .I1(w2), .I2(w3), .I3(w20), .I4(w20), .I5(w20), .I6(w9), .I7(w13), .I8(w20), .I9(w20), .I10(w20), .I11(w20), .I12(w20), .I13(w20), .I14(w20), .I15(w20), .S(ALU_OP), .Z(Result));   //: @(1071,348) /sn:0 /R:1 /w:[ 0 0 0 45 43 39 3 5 35 31 27 23 19 15 11 7 0 0 ] /ss:1 /do:1
  //: joint g35 (w20) @(901, 468) /w:[ 17 18 20 -1 ]
  tran g22(.Z(w11), .I(w9[31]));   //: @(691,545) /sn:0 /R:2 /w:[ 0 1 2 ] /ss:1
  //: joint g31 (w20) @(966, 607) /w:[ 2 4 1 -1 ]
  //: joint g45 (A) @(361, 346) /w:[ 10 9 -1 12 ]
  //: joint g33 (w20) @(938, 468) /w:[ 9 10 12 -1 ]
  //: joint g36 (w20) @(880, 468) /w:[ 21 22 24 -1 ]
  //: joint g41 (w20) @(768, 468) /w:[ 41 42 44 -1 ]
  led g42 (.I(B));   //: @(131,146) /sn:0 /w:[ 7 ] /type:3
  //: joint g40 (w20) @(792, 468) /w:[ 37 38 40 -1 ]
  //: input g12 (ALU_OP) @(1005,123) /sn:0 /w:[ 1 ]
  led g46 (.I(w3));   //: @(681,687) /sn:0 /w:[ 5 ] /type:3
  //: comment g28 /dolink:0 /link:"" @(845,478) /sn:0
  //: /line:"not used pins"
  //: /line:""
  //: /end
  //: joint g34 (w20) @(920, 468) /w:[ 13 14 16 -1 ]
  and g5 (.I0(A), .I1(B), .Z(w1));   //: @(582,191) /sn:0 /w:[ 7 0 1 ]
  //: switch g11 (w23) @(520,372) /sn:0 /w:[ 0 ] /st:0
  //: joint g14 (A) @(361, 322) /w:[ -1 2 1 8 ]
  led g19 (.I(w16));   //: @(610,619) /sn:0 /w:[ 1 ] /type:0
  mux g21 (.I0(w20), .I1(w6), .S(w11), .Z(w13));   //: @(1011,545) /sn:0 /R:2 /w:[ 3 1 1 0 ] /ss:1 /do:1
  //: joint g32 (w20) @(954, 468) /w:[ 5 6 8 -1 ]
  led g20 (.I(w21));   //: @(600,481) /sn:0 /w:[ 1 ] /type:0
  //: joint g43 (B) @(270, 360) /w:[ -1 5 6 8 ]
  Ca2 g0 (.in(B), .out(w0));   //: @(447, 577) /sz:(72, 40) /sn:0 /p:[ Li0>17 Ro0<0 ]
  //: joint g15 (A) @(361, 424) /w:[ 14 13 -1 16 ]
  //: joint g38 (w20) @(836, 468) /w:[ 29 30 32 -1 ]
  //: joint g27 (w13) @(1011, 501) /w:[ 2 4 -1 1 ]
  //: joint g37 (w20) @(862, 468) /w:[ 25 26 28 -1 ]
  //: joint g13 (A) @(361, 277) /w:[ 4 6 -1 3 ]

endmodule

module main;    //: root_module
wire [31:0] w6;    //: /sn:0 {0}(430,382)(527,382){1}
wire w4;    //: /sn:0 {0}(788,317)(673,317){1}
wire [31:0] w3;    //: /sn:0 {0}(673,376)(745,376){1}
wire [31:0] w2;    //: /sn:0 /dp:1 {0}(432,325)(527,325){1}
wire [3:0] w5;    //: /sn:0 /dp:1 {0}(597,226)(597,253)(596,253)(596,281){1}
//: enddecls

  //: dip g4 (w2) @(394,325) /sn:0 /R:1 /w:[ 0 ] /st:0
  led g3 (.I(w3));   //: @(752,376) /sn:0 /R:3 /w:[ 1 ] /type:3
  led g2 (.I(w4));   //: @(795,317) /sn:0 /R:3 /w:[ 0 ] /type:3
  //: dip g1 (w5) @(597,216) /sn:0 /w:[ 0 ] /st:6
  //: dip g5 (w6) @(392,382) /sn:0 /R:1 /w:[ 0 ] /st:0
  ALU g0 (.ALU_OP(w5), .B(w6), .A(w2), .Result(w3), .Zero(w4));   //: @(528, 282) /sz:(144, 125) /sn:0 /p:[ Ti0>1 Li0>1 Li1>1 Ro0<0 Ro1<1 ]

endmodule
