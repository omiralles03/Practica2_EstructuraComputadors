//: version "1.8.7"

module JUMP(PCSrc, SignExtOut, PCNext, Jump, lnm26, PCin);
//: interface  /sz:(118, 106) /bd:[ Ti0>Jump(63/118) Li0>lnm26[25:0](27/106) Li1>PCNext[31:0](57/106) Li2>SignExtOut[31:0](91/106) Bi0>PCSrc(90/118) Ro0<PCin[31:0](52/106) ]
input PCSrc;    //: /sn:0 {0}(510,370)(536,370)(536,311){1}
supply0 w0;    //: /sn:0 {0}(452,261)(452,253)(435,253)(435,274){1}
output [31:0] PCin;    //: /sn:0 /dp:1 {0}(688,278)(626,278){1}
input [31:0] SignExtOut;    //: /sn:0 {0}(361,314)(421,314){1}
input [31:0] PCNext;    //: /sn:0 {0}(286,259)(337,259)(337,282)(370,282){1}
//: {2}(371,282)(403,282){3}
//: {4}(407,282)(421,282){5}
//: {6}(405,280)(405,233)(501,233)(501,278)(520,278){7}
input [25:0] lnm26;    //: /sn:0 /dp:1 {0}(509,217)(343,217){1}
input Jump;    //: /sn:0 {0}(599,342)(613,342)(613,301){1}
wire [5:0] w6;    //: /sn:0 {0}(371,277)(371,207)(509,207){1}
wire [31:0] w7;    //: /sn:0 {0}(515,212)(581,212)(581,268)(597,268){1}
wire w4;    //: /sn:0 {0}(435,322)(435,337)(449,337){1}
wire [31:0] w12;    //: /sn:0 {0}(549,288)(597,288){1}
wire [31:0] w2;    //: /sn:0 {0}(450,298)(520,298){1}
//: enddecls

  //: input g8 (PCSrc) @(508,370) /sn:0 /w:[ 0 ]
  mux g4 (.I0(w12), .I1(w7), .S(Jump), .Z(PCin));   //: @(613,278) /sn:0 /R:1 /w:[ 1 1 1 1 ] /ss:0 /do:0
  add g3 (.A(SignExtOut), .B(PCNext), .S(w2), .CI(w0), .CO(w4));   //: @(437,298) /sn:0 /R:1 /w:[ 1 5 0 1 0 ]
  //: input g2 (SignExtOut) @(359,314) /sn:0 /w:[ 0 ]
  //: input g1 (PCNext) @(284,259) /sn:0 /w:[ 0 ]
  concat g10 (.I0(lnm26), .I1(w6), .Z(w7));   //: @(514,212) /sn:0 /w:[ 0 1 0 ] /dr:0
  //: supply0 g6 (w0) @(452,267) /sn:0 /w:[ 0 ]
  //: joint g9 (PCNext) @(405, 282) /w:[ 4 6 3 -1 ]
  led g7 (.I(w4));   //: @(456,337) /sn:0 /R:3 /w:[ 1 ] /type:0
  //: input g12 (Jump) @(597,342) /sn:0 /w:[ 0 ]
  tran g11(.Z(w6), .I(PCNext[31:26]));   //: @(371,280) /sn:0 /R:1 /w:[ 0 1 2 ] /ss:0
  mux g5 (.I0(PCNext), .I1(w2), .S(PCSrc), .Z(w12));   //: @(536,288) /sn:0 /R:1 /w:[ 7 1 1 0 ] /ss:0 /do:1
  //: input g0 (lnm26) @(341,217) /sn:0 /w:[ 1 ]
  //: output g13 (PCin) @(685,278) /sn:0 /w:[ 0 ]

endmodule

module MEM(WriteData, ReadData, MemWrite, MemRead, Address);
//: interface  /sz:(130, 124) /bd:[ Ti0>MemWrite(56/130) Li0>Address[31:0](31/124) Li1>WriteData[31:0](101/124) Bi0>MemRead(64/130) Ro0<ReadData[31:0](44/124) ]
output [31:0] ReadData;    //: /sn:0 {0}(644,286)(644,315){1}
//: {2}(646,317)(690,317){3}
//: {4}(642,317)(607,317){5}
input [31:0] WriteData;    //: /sn:0 /dp:1 {0}(607,235)(644,235)(644,270){1}
input MemWrite;    //: /sn:0 {0}(567,271)(588,271){1}
//: {2}(592,271)(606,271)(606,262)(662,262)(662,278)(649,278){3}
//: {4}(590,273)(590,294){5}
input MemRead;    //: /sn:0 {0}(631,373)(597,373)(597,344){1}
supply0 w5;    //: /sn:0 {0}(583,371)(583,344){1}
input [31:0] Address;    //: /sn:0 {0}(512,319)(572,319){1}
//: enddecls

  bufif1 g8 (.Z(ReadData), .I(WriteData), .E(MemWrite));   //: @(644,276) /sn:0 /R:3 /w:[ 0 1 3 ]
  //: input g4 (WriteData) @(605,235) /sn:0 /w:[ 0 ]
  //: output g3 (ReadData) @(687,317) /sn:0 /w:[ 3 ]
  //: input g2 (MemWrite) @(565,271) /sn:0 /w:[ 0 ]
  //: input g1 (MemRead) @(633,373) /sn:0 /R:2 /w:[ 0 ]
  //: joint g10 (ReadData) @(644, 317) /w:[ 2 1 4 -1 ]
  //: supply0 g6 (w5) @(583,377) /sn:0 /w:[ 0 ]
  //: joint g9 (MemWrite) @(590, 271) /w:[ 2 -1 1 4 ]
  //: comment g7 /dolink:0 /link:"" @(396,417) /sn:0
  //: /line:"lw: (CS & WE) = 0, MemWrite 1, valor de @Adress surt per ReadData"
  //: /line:"sw: (CS & OE) = 0, WriteData 1, guarda valor WriteData a @Adress"
  //: /end
  ram g5 (.A(Address), .D(ReadData), .WE(MemWrite), .OE(MemRead), .CS(w5));   //: @(590,318) /sn:0 /w:[ 1 5 5 1 1 ]
  //: input g0 (Address) @(510,319) /sn:0 /w:[ 0 ]

endmodule

module Zero(f, i);
//: interface  /sz:(40, 40) /bd:[ Li0>i[31:0](21/40) Li1>i[31:0](21/40) Li2>i[31:0](21/40) Ro0<f(22/40) Ro1<f(22/40) Ro2<f(22/40) ]
supply0 w0;    //: /sn:0 {0}(803,314)(803,304)(788,304)(788,362)(779,362)(779,372){1}
input f;    //: /sn:0 {0}(769,401)(769,481)(804,481)(804,441)(873,441)(873,448)(929,448)(929,393)(899,393){1}
input [31:0] i;    //: /sn:0 {0}(276,291)(433,291)(433,299)(443,299){1}
supply1 w2;    //: /sn:0 {0}(750,325)(750,368)(759,368)(759,372){1}
wire [31:0] w7;    //: /sn:0 {0}(517,298)(575,298)(575,302)(676,302){1}
//: {2}(677,302)(713,302)(713,268)(787,268)(787,239){3}
wire [31:0] w1;    //: /sn:0 /dp:1 {0}(496,228)(496,252)(574,252){1}
wire o;    //: /sn:0 {0}(677,306)(677,327){1}
//: {2}(675,329)(600,329)(600,402)(615,402)(615,392){3}
//: {4}(677,331)(677,388)(746,388){5}
//: enddecls

  led g4 (.I(w7));   //: @(787,232) /sn:0 /w:[ 3 ] /type:3
  //: joint g8 (o) @(677, 329) /w:[ -1 1 2 4 ]
  //: dip g3 (w1) @(496,218) /sn:0 /w:[ 0 ] /st:0
  Ca2 g2 (.in(i), .out(w7));   //: @(444, 277) /sz:(72, 40) /sn:0 /p:[ Li0>1 Ro0<0 ]
  //: input g1 (f) @(897,393) /sn:0 /w:[ 1 ]
  //: supply0 g10 (w0) @(803,320) /sn:0 /w:[ 0 ]
  mux g6 (.I0(w2), .I1(w0), .S(o), .Z(f));   //: @(769,388) /sn:0 /w:[ 1 1 5 0 ] /ss:0 /do:0
  led g7 (.I(o));   //: @(615,385) /sn:0 /w:[ 3 ] /type:0
  //: supply1 g9 (w2) @(761,325) /sn:0 /w:[ 0 ]
  tran g5(.Z(o), .I(w7[31]));   //: @(677,300) /sn:0 /R:1 /w:[ 0 1 2 ] /ss:1
  //: input g0 (i) @(274,291) /sn:0 /w:[ 0 ]

endmodule

module READ(clk, Read2, RegWrite, Read1, WriteData, RegDst, Write, SignExtIn, clr, Data1, Data2, SignExtOut);
//: interface  /sz:(173, 238) /bd:[ Ti0>RegWrite(85/173) Li0>Read1[4:0](29/238) Li1>Read2[4:0](70/238) Li2>Write[4:0](106/238) Li3>WriteData[31:0](174/238) Li4>SignExtIn[15:0](205/238) Li5>RegDst(140/238) Bi0>clk(57/173) Bi1>clr(119/173) Ro0<SignExtOut[31:0](208/238) Ro1<Data2[31:0](140/238) Ro2<Data1[31:0](78/238) ]
output [31:0] Data2;    //: /sn:0 {0}(689,234)(621,234){1}
input [4:0] Write;    //: {0}(336,213)(388,213){1}
input [31:0] WriteData;    //: /sn:0 {0}(389,296)(441,296)(441,243)(472,243){1}
output [31:0] SignExtOut;    //: /sn:0 /dp:1 {0}(722,399)(654,399){1}
output [31:0] Data1;    //: /sn:0 /dp:1 {0}(695,142)(621,142){1}
input RegDst;    //: /sn:0 {0}(333,252)(404,252)(404,226){1}
input RegWrite;    //: /sn:0 {0}(513,310)(513,278){1}
input clr;    //: /sn:0 {0}(506,74)(539,74)(539,94){1}
input clk;    //: /sn:0 {0}(581,306)(581,278){1}
input [4:0] Read1;    //: /sn:0 {0}(364,127)(472,127){1}
input [4:0] Read2;    //: /sn:0 /dp:1 {0}(329,167)(361,167){1}
//: {2}(365,167)(472,167){3}
//: {4}(363,169)(363,193)(388,193){5}
input [15:0] SignExtIn;    //: /sn:0 /dp:1 {0}(352,400)(445,400){1}
wire [4:0] w6;    //: /sn:0 /dp:1 {0}(417,203)(472,203){1}
//: enddecls

  //: input g4 (clk) @(581,308) /sn:0 /R:1 /w:[ 0 ]
  //: input g8 (Read2) @(327,167) /sn:0 /w:[ 0 ]
  //: input g3 (RegWrite) @(513,312) /sn:0 /R:1 /w:[ 0 ]
  //: input g2 (Read1) @(362,127) /sn:0 /w:[ 0 ]
  SignExtend g1 (.lnm16(SignExtIn), .D32b(SignExtOut));   //: @(446, 363) /sz:(207, 73) /sn:0 /p:[ Li0>1 Ro0<1 ]
  //: input g10 (WriteData) @(387,296) /sn:0 /w:[ 0 ]
  mux g6 (.I0(Read2), .I1(Write), .S(RegDst), .Z(w6));   //: @(404,203) /sn:0 /R:1 /w:[ 5 1 1 0 ] /ss:0 /do:1
  //: input g7 (RegDst) @(331,252) /sn:0 /w:[ 0 ]
  //: input g9 (Write) @(334,213) /sn:0 /w:[ 0 ]
  //: input g12 (SignExtIn) @(350,400) /sn:0 /w:[ 0 ]
  //: input g5 (clr) @(504,74) /sn:0 /w:[ 0 ]
  //: joint g11 (Read2) @(363, 167) /w:[ 2 -1 1 4 ]
  //: output g14 (Data1) @(692,142) /sn:0 /w:[ 0 ]
  BRegs32x32 g0 (.clr(clr), .Read1(Read1), .Read2(Read2), .Write(w6), .WriteData(WriteData), .clk(clk), .RegWrite(RegWrite), .Data1(Data1), .Data2(Data2));   //: @(473, 95) /sz:(147, 182) /sn:0 /p:[ Ti0>1 Li0>1 Li1>3 Li2>1 Li3>1 Bi0>1 Bi1>1 Ro0<1 Ro1<1 ]
  //: output g15 (Data2) @(686,234) /sn:0 /w:[ 0 ]
  //: output g13 (SignExtOut) @(719,399) /sn:0 /w:[ 0 ]

endmodule

module SignExtend(D32b, lnm16);
//: interface  /sz:(207, 73) /bd:[ Li0>lnm16[15:0](37/73) Ro0<D32b[31:0](36/73) ]
output [31:0] D32b;    //: /sn:0 /dp:1 {0}(513,367)(476,367){1}
input [15:0] lnm16;    //: /sn:0 /dp:3 {0}(470,372)(388,372)(388,413)(350,413){1}
//: {2}(349,413)(188,413){3}
wire [15:0] w6;    //: /sn:0 /dp:1 {0}(270,298)(302,298)(302,280)(334,280){1}
wire w4;    //: /sn:0 {0}(350,408)(350,293){1}
wire [15:0] w0;    //: /sn:0 /dp:1 {0}(270,244)(303,244)(303,260)(334,260){1}
wire [15:0] w1;    //: /sn:0 /dp:1 {0}(470,362)(388,362)(388,270)(363,270){1}
//: enddecls

  //: dip g4 (w6) @(232,298) /sn:0 /R:1 /w:[ 0 ] /st:0
  //: comment g8 /dolink:0 /link:"" @(188,321) /sn:0 /R:1
  //: /line:"0xb0000000000000000"
  //: /end
  //: output g3 (D32b) @(510,367) /sn:0 /w:[ 0 ]
  concat g2 (.I0(lnm16), .I1(w1), .Z(D32b));   //: @(475,367) /sn:0 /w:[ 0 0 1 ] /dr:0
  mux g1 (.I0(w6), .I1(w0), .S(w4), .Z(w1));   //: @(350,270) /sn:0 /R:1 /w:[ 1 1 1 1 ] /ss:0 /do:0
  tran g6(.Z(w4), .I(lnm16[15]));   //: @(350,411) /sn:0 /R:1 /w:[ 0 2 1 ] /ss:0
  //: comment g7 /dolink:0 /link:"" @(189,200) /sn:0 /R:1
  //: /line:"0xb1111111111111111"
  //: /end
  //: comment g9 /dolink:0 /link:"" @(222,180) /sn:0 /R:1
  //: /line:"65535"
  //: /end
  //: dip g5 (w0) @(232,244) /sn:0 /R:1 /w:[ 0 ] /st:65535
  //: input g0 (lnm16) @(186,413) /sn:0 /w:[ 3 ]

endmodule

module DataMemory(ReadData, MemWrite, MemRead, WriteData, Address);
//: interface  /sz:(113, 152) /bd:[ Ti0>MemWrite(49/113) Li0>Address[31:0](39/152) Li1>WriteData[31:0](125/152) Bi0>MemRead(56/113) Ro0<ReadData[31:0](54/152) Ro1<DataMemory[31:0](105/152) ]
output [31:0] ReadData;    //: /sn:0 /dp:1 {0}(479,279)(628,279)(628,363){1}
//: {2}(630,365)(714,365)(714,391)(829,391){3}
//: {4}(626,365)(586,365){5}
input [31:0] WriteData;    //: /sn:0 {0}(463,279)(423,279)(423,241)(128,241){1}
input MemWrite;    //: /sn:0 /dp:1 {0}(569,342)(569,333)(230,333){1}
//: {2}(228,331)(228,178)(471,178)(471,274){3}
//: {4}(228,335)(228,436)(198,436){5}
//: {6}(194,436)(134,436)(134,375)(64,375){7}
//: {8}(196,438)(196,471)(281,471){9}
input MemRead;    //: /sn:0 {0}(576,392)(576,567)(225,567)(225,509){1}
//: {2}(227,507)(273,507)(273,476)(281,476){3}
//: {4}(223,507)(49,507){5}
input [31:0] Address;    //: /sn:0 {0}(336,367)(551,367){1}
wire w0;    //: /sn:0 {0}(562,392)(562,474)(302,474){1}
//: enddecls

  ram g4 (.A(Address), .D(ReadData), .WE(!MemWrite), .OE(!MemRead), .CS(w0));   //: @(569,366) /sn:0 /w:[ 1 5 0 0 0 ]
  //: output g8 (ReadData) @(826,391) /sn:0 /w:[ 3 ]
  //: comment g3 /dolink:0 /link:"" @(199,90) /sn:0
  //: /line:"case1: lw Memread=1 MemWrite=0 MTR=1"
  //: /line:"case2: sw Memread=0 MemWrite=1 MTR=X"
  //: /end
  //: input g2 (MemWrite) @(62,375) /sn:0 /w:[ 7 ]
  //: comment g1 /dolink:0 /link:"" @(293,493) /sn:0
  //: /line:"Mr   Mw"
  //: /line:"0    0    1"
  //: /line:"0    1    0"
  //: /line:"1    0    0"
  //: /line:"1    1    1"
  //: /end
  //: input g10 (MemRead) @(47,507) /sn:0 /w:[ 5 ]
  bufif1 g6 (.Z(ReadData), .I(WriteData), .E(MemWrite));   //: @(469,279) /sn:0 /w:[ 0 0 3 ]
  xnor g9 (.I0(MemWrite), .I1(MemRead), .Z(w0));   //: @(292,474) /sn:0 /w:[ 9 3 1 ]
  //: input g7 (WriteData) @(126,241) /sn:0 /w:[ 1 ]
  //: joint g12 (MemWrite) @(196, 436) /w:[ 5 -1 6 8 ]
  //: joint g14 (MemRead) @(225, 507) /w:[ 2 -1 4 1 ]
  //: input g5 (Address) @(334,367) /sn:0 /w:[ 0 ]
  //: joint g11 (ReadData) @(628, 365) /w:[ 2 1 4 -1 ]
  //: comment g0 /dolink:0 /link:"" @(615,414) /sn:0
  //: /line:"lw: if (CS & OE) = 0, valor dins @Adress surt per D"
  //: /line:"sw: if (CS & WE) = 0, D es guarda a @Adress"
  //: /line:""
  //: /end
  //: joint g13 (MemWrite) @(228, 333) /w:[ 1 2 -1 4 ]

endmodule

module ALU(Result, Zero, B, A, ALU_OP);
//: interface  /sz:(94, 87) /bd:[ Ti0>ALU_OP[3:0](45/94) Ti1>ALU_OP[3:0](45/94) Ti2>ALU_OP[3:0](45/94) Ti3>ALU_OP[3:0](45/94) Li0>A[31:0](30/87) Li1>B[31:0](70/87) Li2>B[31:0](70/87) Li3>A[31:0](30/87) Li4>A[31:0](30/87) Li5>B[31:0](70/87) Li6>B[31:0](70/87) Li7>A[31:0](30/87) Ro0<Zero(32/87) Ro1<Result[31:0](66/87) Ro2<Result[31:0](66/87) Ro3<Zero(32/87) Ro4<Zero(32/87) Ro5<Result[31:0](66/87) Ro6<Result[31:0](66/87) Ro7<Zero(32/87) ]
input [31:0] B;    //: /sn:0 /dp:1 {0}(571,193)(270,193)(270,280){1}
//: {2}(272,282)(576,282){3}
//: {4}(270,284)(270,358){5}
//: {6}(268,360)(131,360)(131,153){7}
//: {8}(270,362)(270,411){9}
//: {10}(268,413)(222,413){11}
//: {12}(270,415)(270,454){13}
//: {14}(272,456)(569,456){15}
//: {16}(270,458)(270,599)(446,599){17}
output Zero;    //: /sn:0 {0}(1411,566)(1505,566){1}
input [31:0] A;    //: /sn:0 {0}(317,322)(359,322){1}
//: {2}(361,320)(361,279){3}
//: {4}(363,277)(576,277){5}
//: {6}(361,275)(361,188)(571,188){7}
//: {8}(361,324)(361,344){9}
//: {10}(363,346)(513,346)(513,112){11}
//: {12}(361,348)(361,422){13}
//: {14}(363,424)(569,424){15}
//: {16}(361,426)(361,566)(570,566){17}
output [31:0] Result;    //: /sn:0 /dp:1 {0}(1098,341)(1317,341){1}
//: {2}(1321,341)(1415,341){3}
//: {4}(1319,343)(1319,565)(1369,565){5}
supply0 [31:0] w1;    //: /sn:0 /dp:2 {0}(1069,337)(932,337)(932,342){1}
//: {2}(934,344)(1069,344){3}
//: {4}(932,346)(932,348){5}
//: {6}(934,350)(1069,350){7}
//: {8}(932,352)(932,419){9}
input [3:0] ALU_OP;    //: /sn:0 /dp:3 {0}(1025,129)(995,129){1}
//: {2}(994,129)(929,129){3}
wire [31:0] w6;    //: /sn:0 /dp:1 {0}(1021,699)(1021,561){1}
wire [31:0] w13;    //: /sn:0 {0}(1011,532)(1011,503){1}
//: {2}(1013,501)(1162,501)(1162,493){3}
//: {4}(1011,499)(1011,364)(1069,364){5}
wire w16;    //: /sn:0 {0}(584,606)(584,636)(610,636)(610,626){1}
wire [2:0] w7;    //: /sn:0 {0}(995,133)(995,268)(1085,268)(1085,318){1}
wire [31:0] w4;    //: /sn:0 {0}(1069,317)(1043,317)(1043,304)(704,304)(704,191)(592,191){1}
wire [31:0] w3;    //: /sn:0 /dp:1 {0}(685,683)(685,643)(676,643)(676,584){1}
//: {2}(678,582)(693,582)(693,545){3}
//: {4}(693,544)(693,357)(1069,357){5}
//: {6}(674,582)(599,582){7}
wire w22;    //: /sn:0 {0}(545,525)(584,525)(584,558){1}
wire [31:0] w0;    //: /sn:0 {0}(520,598)(570,598){1}
wire [31:0] w20;    //: /sn:0 {0}(953,644)(953,607)(1001,607)(1001,561){1}
wire w23;    //: /sn:0 {0}(537,372)(583,372)(583,416){1}
wire w21;    //: /sn:0 {0}(583,464)(583,498)(600,498)(600,488){1}
wire w11;    //: /sn:0 {0}(697,545)(988,545){1}
wire [31:0] w2;    //: /sn:0 {0}(597,280)(693,280)(693,324)(1069,324){1}
wire [31:0] w5;    //: /sn:0 {0}(598,440)(656,440)(656,330)(1069,330){1}
//: enddecls

  add g8 (.A(w0), .B(A), .S(w3), .CI(w22), .CO(w16));   //: @(586,582) /sn:0 /R:1 /w:[ 1 17 7 1 0 ]
  //: output g4 (Result) @(1412,341) /sn:0 /w:[ 3 ]
  led g44 (.I(A));   //: @(513,105) /sn:0 /w:[ 11 ] /type:3
  //: joint g16 (B) @(270, 282) /w:[ 2 1 -1 4 ]
  //: output g3 (Zero) @(1502,566) /sn:0 /w:[ 1 ]
  led g26 (.I(w13));   //: @(1162,486) /sn:0 /w:[ 3 ] /type:3
  //: joint g17 (B) @(270, 413) /w:[ -1 9 10 12 ]
  //: input g2 (B) @(220,413) /sn:0 /w:[ 11 ]
  //: comment g23 /dolink:0 /link:"" @(1052,527) /sn:0
  //: /line:"if (A < B)   // bit 31 = 1"
  //: /line:"   ALU = 1;"
  //: /line:"else         // bit 31 = 0"
  //: /line:"   ALU = 0;"
  //: /end
  //: joint g30 (w13) @(1011, 501) /w:[ 2 4 -1 1 ]
  //: dip g24 (w6) @(1021,710) /sn:0 /R:2 /w:[ 0 ] /st:1
  //: input g1 (A) @(315,322) /sn:0 /w:[ 0 ]
  Zero g29 (.i(Result), .f(Zero));   //: @(1370, 544) /sz:(40, 40) /sn:0 /p:[ Li0>5 Ro0<0 ]
  //: joint g18 (B) @(270, 456) /w:[ 14 13 -1 16 ]
  //: dip g25 (w20) @(953,655) /sn:0 /R:2 /w:[ 0 ] /st:0
  //: switch g10 (w22) @(528,525) /sn:0 /w:[ 0 ] /st:0
  or g6 (.I0(A), .I1(B), .Z(w2));   //: @(587,280) /sn:0 /w:[ 5 3 0 ]
  add g9 (.A(B), .B(A), .S(w5), .CI(w23), .CO(w21));   //: @(585,440) /sn:0 /R:1 /w:[ 15 15 0 1 0 ]
  mux g7 (.I0(w4), .I1(w2), .I2(w5), .I3(w1), .I4(w1), .I5(w1), .I6(w3), .I7(w13), .S(w7), .Z(Result));   //: @(1085,341) /sn:0 /R:1 /w:[ 0 1 1 0 3 7 5 5 1 0 ] /ss:1 /do:1
  //: joint g35 (Result) @(1319, 341) /w:[ 2 -1 1 4 ]
  tran g22(.Z(w11), .I(w3[31]));   //: @(691,545) /sn:0 /R:2 /w:[ 0 3 4 ] /ss:1
  //: joint g31 (w3) @(676, 582) /w:[ 2 -1 6 1 ]
  //: joint g45 (A) @(361, 346) /w:[ 10 9 -1 12 ]
  //: joint g33 (w1) @(932, 344) /w:[ 2 1 -1 4 ]
  led g42 (.I(B));   //: @(131,146) /sn:0 /w:[ 7 ] /type:3
  //: input g12 (ALU_OP) @(927,129) /sn:0 /w:[ 3 ]
  //: comment g28 /dolink:0 /link:"" @(846,413) /sn:0
  //: /line:"not used pins"
  //: /line:""
  //: /end
  led g46 (.I(w3));   //: @(685,690) /sn:0 /R:2 /w:[ 0 ] /type:3
  //: joint g34 (w1) @(932, 350) /w:[ 6 5 -1 8 ]
  //: joint g14 (A) @(361, 322) /w:[ -1 2 1 8 ]
  //: switch g11 (w23) @(520,372) /sn:0 /w:[ 0 ] /st:0
  and g5 (.I0(A), .I1(B), .Z(w4));   //: @(582,191) /sn:0 /w:[ 7 0 1 ]
  mux g21 (.I0(w20), .I1(w6), .S(w11), .Z(w13));   //: @(1011,545) /sn:0 /R:2 /w:[ 1 1 1 0 ] /ss:1 /do:1
  led g19 (.I(w16));   //: @(610,619) /sn:0 /w:[ 1 ] /type:0
  led g20 (.I(w21));   //: @(600,481) /sn:0 /w:[ 1 ] /type:0
  //: supply0 g32 (w1) @(932,425) /sn:0 /w:[ 9 ]
  //: joint g15 (A) @(361, 424) /w:[ 14 13 -1 16 ]
  Ca2 g0 (.in(B), .out(w0));   //: @(447, 577) /sz:(72, 40) /sn:0 /p:[ Li0>17 Ro0<0 ]
  //: joint g43 (B) @(270, 360) /w:[ -1 5 6 8 ]
  tran g27(.Z(w7), .I(ALU_OP[2:0]));   //: @(995,127) /sn:0 /R:1 /w:[ 0 2 1 ] /ss:1
  //: joint g13 (A) @(361, 277) /w:[ 4 6 -1 3 ]

endmodule

module EXE(Zero, Result, ALU_OP, B, A);
//: interface  /sz:(160, 125) /bd:[ Ti0>ALU_OP[3:0](79/160) Li0>A[31:0](51/125) Li1>B[31:0](96/125) Ro0<Result[31:0](86/125) Ro1<Zero(48/125) ]
input [31:0] B;    //: /sn:0 {0}(349,318)(396,318){1}
//: {2}(398,316)(398,297){3}
//: {4}(400,295)(530,295){5}
//: {6}(398,293)(398,212){7}
//: {8}(400,210)(524,210){9}
//: {10}(398,208)(398,162)(523,162){11}
//: {12}(398,320)(398,530)(444,530){13}
output Zero;    //: /sn:0 /dp:1 {0}(860,324)(896,324){1}
supply0 w3;    //: /sn:0 {0}(439,464)(439,453)(458,453)(458,490){1}
supply0 w0;    //: /sn:0 {0}(528,239)(528,224)(544,224)(544,255){1}
input [31:0] A;    //: /sn:0 /dp:1 {0}(523,157)(444,157)(444,203){1}
//: {2}(446,205)(524,205){3}
//: {4}(444,207)(444,261){5}
//: {6}(446,263)(530,263){7}
//: {8}(442,263)(352,263){9}
//: {10}(444,265)(444,429)(536,429){11}
output [31:0] Result;    //: /sn:0 {0}(886,290)(807,290){1}
//: {2}(803,290)(791,290){3}
//: {4}(805,292)(805,324)(839,324){5}
input [3:0] ALU_OP;    //: /sn:0 {0}(740,204)(777,204){1}
//: {2}(778,204)(784,204){3}
supply0 w26;    //: /sn:0 {0}(536,400)(536,390)(550,390)(550,421){1}
wire [31:0] w6;    //: /sn:0 /dp:1 {0}(762,273)(665,273)(665,208)(545,208){1}
wire [31:0] w13;    //: /sn:0 /dp:3 {0}(565,445)(645,445)(645,437){1}
//: {2}(645,436)(645,376)(702,376)(702,306)(762,306){3}
wire [2:0] w7;    //: /sn:0 {0}(778,208)(778,267){1}
wire [31:0] w4;    //: /sn:0 /dp:1 {0}(762,266)(683,266)(683,160)(544,160){1}
wire w25;    //: /sn:0 {0}(544,303)(544,331){1}
wire [31:0] w20;    //: /sn:0 {0}(689,494)(689,474){1}
//: {2}(691,472)(727,472)(727,453){3}
//: {4}(689,470)(689,293)(699,293){5}
//: {6}(703,293)(762,293){7}
//: {8}(701,291)(701,286)(762,286){9}
//: {10}(701,295)(701,299)(762,299){11}
wire [31:0] w19;    //: /sn:0 /dp:1 {0}(737,424)(737,313)(762,313){1}
wire w10;    //: /sn:0 {0}(458,538)(458,560){1}
wire [31:0] w1;    //: /sn:0 /dp:1 {0}(353,498)(444,498){1}
wire [31:0] w8;    //: /sn:0 {0}(473,514)(513,514)(513,461)(536,461){1}
wire w17;    //: /sn:0 {0}(649,437)(714,437){1}
wire w14;    //: /sn:0 /dp:1 {0}(550,489)(550,469){1}
wire [31:0] w11;    //: /sn:0 /dp:1 {0}(762,279)(559,279){1}
wire [31:0] w5;    //: /sn:0 /dp:1 {0}(747,453)(747,473)(786,473)(786,493){1}
//: enddecls

  add g8 (.A(w8), .B(A), .S(w13), .CI(w26), .CO(w14));   //: @(552,445) /sn:0 /R:1 /w:[ 1 11 0 1 1 ]
  //: output g4 (Zero) @(893,324) /sn:0 /w:[ 1 ]
  led g16 (.I(w25));   //: @(544,338) /sn:0 /R:2 /w:[ 1 ] /type:3
  //: output g3 (Result) @(883,290) /sn:0 /w:[ 0 ]
  //: dip g26 (w20) @(689,505) /sn:0 /R:2 /w:[ 0 ] /st:0
  //: joint g17 (A) @(444, 263) /w:[ 6 5 8 10 ]
  //: input g2 (ALU_OP) @(738,204) /sn:0 /w:[ 0 ]
  //: comment g30 /dolink:0 /link:"" @(597,289) /sn:0 /R:2
  //: /line:"not used pins"
  //: /line:"    0011"
  //: /line:"    0100"
  //: /line:"    0101"
  //: /line:"   "
  //: /end
  mux g23 (.I0(w4), .I1(w6), .I2(w11), .I3(w20), .I4(w20), .I5(w20), .I6(w13), .I7(w19), .S(w7), .Z(Result));   //: @(778,290) /sn:0 /R:1 /w:[ 0 0 0 9 7 11 3 1 1 3 ] /ss:1 /do:1
  mux g24 (.I0(w20), .I1(w5), .S(w17), .Z(w19));   //: @(737,437) /sn:0 /R:2 /w:[ 3 0 1 0 ] /ss:1 /do:1
  //: input g1 (B) @(347,318) /sn:0 /w:[ 0 ]
  //: joint g29 (w20) @(701, 293) /w:[ 6 8 5 10 ]
  //: joint g18 (B) @(398, 210) /w:[ 8 10 -1 7 ]
  tran g25(.Z(w17), .I(w13[31]));   //: @(643,437) /sn:0 /R:2 /w:[ 0 1 2 ] /ss:1
  add g10 (.A(B), .B(A), .S(w11), .CI(w0), .CO(w25));   //: @(546,279) /sn:0 /R:1 /w:[ 5 7 1 1 0 ]
  or g6 (.I0(A), .I1(B), .Z(w6));   //: @(535,208) /sn:0 /w:[ 3 9 1 ]
  led g9 (.I(w10));   //: @(458,567) /sn:0 /R:2 /w:[ 1 ] /type:3
  add g7 (.A(!B), .B(w1), .S(w8), .CI(w3), .CO(w10));   //: @(460,514) /sn:0 /R:1 /w:[ 13 1 0 1 0 ]
  tran g31(.Z(w7), .I(ALU_OP[2:0]));   //: @(778,202) /sn:0 /R:1 /w:[ 0 1 2 ] /ss:1
  //: comment g22 /dolink:0 /link:"" @(481,522) /sn:0 /R:1
  //: /line:"Ca2"
  //: /end
  //: joint g33 (Result) @(805, 290) /w:[ 1 -1 2 4 ]
  //: supply0 g12 (w0) @(528,245) /sn:0 /w:[ 0 ]
  //: comment g34 /dolink:0 /link:"" @(614,536) /sn:0 /R:2
  //: /line:"A <  B -> b31 = 1 -> Result = 1"
  //: /line:"A >= B -> b31 = 0 -> Result = 0"
  //: /line:"    "
  //: /end
  //: joint g28 (w20) @(689, 472) /w:[ 2 4 -1 1 ]
  //: supply0 g14 (w26) @(536,406) /sn:0 /w:[ 0 ]
  //: joint g11 (A) @(444, 205) /w:[ 2 1 -1 4 ]
  and g5 (.I0(A), .I1(B), .Z(w4));   //: @(534,160) /sn:0 /w:[ 0 11 1 ]
  //: dip g21 (w1) @(315,498) /sn:0 /R:1 /w:[ 0 ] /st:1
  //: joint g19 (B) @(398, 295) /w:[ 4 6 -1 3 ]
  nor g32 (.I0(Result), .Z(Zero));   //: @(850,324) /sn:0 /w:[ 5 0 ]
  //: joint g20 (B) @(398, 318) /w:[ -1 2 1 12 ]
  led g15 (.I(w14));   //: @(550,496) /sn:0 /R:2 /w:[ 0 ] /type:3
  //: input g0 (A) @(350,263) /sn:0 /w:[ 9 ]
  //: dip g27 (w5) @(786,504) /sn:0 /R:2 /w:[ 1 ] /st:1
  //: supply0 g13 (w3) @(439,470) /sn:0 /w:[ 0 ]

endmodule

module BRegs32x32(Read2, Write, Read1, Data2, Data1, clr, clk, RegWrite, WriteData);
//: interface  /sz:(147, 182) /bd:[ Ti0>clr(66/147) Li0>Read1[4:0](32/182) Li1>Read2[4:0](72/182) Li2>Write[4:0](108/182) Li3>WriteData[31:0](148/182) Bi0>clk(108/147) Bi1>RegWrite(40/147) Ro0<Data1[31:0](47/182) Ro1<Data2[31:0](139/182) ]
output [31:0] Data2;    //: /sn:0 {0}(668,485)(668,472)(669,472)(669,445){1}
input [4:0] Write;    //: /sn:0 {0}(-238,-38)(-138,-38)(-138,-37)(-66,-37){1}
//: {2}(-65,-37)(-28,-37){3}
//: {4}(-27,-37)(-16,-37){5}
input [31:0] WriteData;    //: /sn:0 {0}(669,157)(669,75)(481,75){1}
//: {2}(477,75)(292,75){3}
//: {4}(288,75)(89,75){5}
//: {6}(85,75)(-104,75)(-104,73)(-237,73){7}
//: {8}(87,77)(87,157){9}
//: {10}(290,77)(290,107)(291,107)(291,152){11}
//: {12}(479,77)(479,157){13}
output [31:0] Data1;    //: /sn:0 {0}(59,382)(59,465){1}
supply1 w21;    //: /sn:0 {0}(82,3)(57,3)(57,-11){1}
input clr;    //: /sn:0 {0}(721,193)(731,193)(731,-83)(543,-83){1}
//: {2}(539,-83)(355,-83){3}
//: {4}(351,-83)(150,-83){5}
//: {6}(146,-83)(-44,-83)(-44,-92)(-235,-92){7}
//: {8}(148,-81)(148,193)(139,193){9}
//: {10}(353,-81)(353,188)(343,188){11}
//: {12}(541,-81)(541,193)(531,193){13}
input RegWrite;    //: /sn:0 {0}(-237,263)(-71,263){1}
//: {2}(-67,263)(171,263){3}
//: {4}(175,263)(370,263){5}
//: {6}(374,263)(552,263)(552,219)(556,219){7}
//: {8}(372,261)(372,219)(383,219){9}
//: {10}(173,261)(173,214)(183,214){11}
//: {12}(-69,261)(-69,219)(-38,219){13}
input clk;    //: /sn:0 {0}(556,214)(542,214)(542,285)(364,285){1}
//: {2}(362,283)(362,214)(383,214){3}
//: {4}(360,285)(167,285){5}
//: {6}(165,283)(165,209)(183,209){7}
//: {8}(163,285)(-56,285){9}
//: {10}(-58,283)(-58,214)(-38,214){11}
//: {12}(-60,285)(-237,285){13}
input [4:0] Read1;    //: {0}(-237,96)(-208,96)(-208,95)(-124,95){1}
//: {2}(-123,95)(-96,95){3}
//: {4}(-95,95)(-78,95){5}
input [4:0] Read2;    //: {0}(-237,145)(-141,145){1}
//: {2}(-140,145)(-123,145)(-123,144)(-94,144){3}
//: {4}(-93,144)(-79,144){5}
wire [1:0] w6;    //: /sn:0 {0}(36,369)(-123,369)(-123,99){1}
wire w16;    //: /sn:0 {0}(39,205)(-50,205)(-50,39)(88,39)(88,19){1}
wire w4;    //: /sn:0 {0}(112,19)(112,46)(370,46)(370,205)(431,205){1}
wire [31:0] w3;    //: /sn:0 {0}(77,353)(77,334)(659,334)(659,228){1}
wire [31:0] R2;    //: {0}(65,353)(65,319)(469,319)(469,228){1}
wire [31:0] w0;    //: /sn:0 {0}(651,416)(651,398)(105,398)(105,228){1}
wire w22;    //: /sn:0 {0}(404,217)(431,217){1}
wire w20;    //: /sn:0 {0}(124,19)(124,29)(556,29)(556,205)(621,205){1}
wire [2:0] w19;    //: /sn:0 {0}(431,169)(419,169)(419,109){1}
//: {2}(421,107)(606,107)(606,169)(621,169){3}
//: {4}(417,107)(297,107)(297,106)(231,106){5}
//: {6}(227,106)(25,106){7}
//: {8}(21,106)(-95,106)(-95,99){9}
//: {10}(23,108)(23,169)(39,169){11}
//: {12}(229,108)(229,164)(243,164){13}
wire [2:0] w18;    //: /sn:0 {0}(431,180)(402,180)(402,125){1}
//: {2}(404,123)(589,123)(589,180)(621,180){3}
//: {4}(400,123)(279,123)(279,122)(212,122){5}
//: {6}(208,122)(8,122){7}
//: {8}(4,122)(-93,122)(-93,139){9}
//: {10}(6,124)(6,180)(39,180){11}
//: {12}(210,124)(210,175)(243,175){13}
wire w23;    //: /sn:0 {0}(577,217)(621,217){1}
wire [1:0] w10;    //: /sn:0 {0}(-140,149)(-140,432)(646,432){1}
wire [2:0] w24;    //: /sn:0 {0}(431,193)(381,193)(381,141){1}
//: {2}(383,139)(568,139)(568,193)(621,193){3}
//: {4}(379,139)(260,139)(260,138)(195,138){5}
//: {6}(191,138)(-13,138){7}
//: {8}(-17,138)(-65,138)(-65,-33){9}
//: {10}(-15,140)(-15,193)(39,193){11}
//: {12}(193,140)(193,188)(243,188){13}
wire w31;    //: /sn:0 {0}(243,200)(178,200)(178,60)(100,60)(100,19){1}
wire w1;    //: /sn:0 {0}(-17,217)(39,217){1}
wire [31:0] R1;    //: {0}(281,223)(281,308)(53,308)(53,353){1}
wire [31:0] R3;    //: {0}(687,228)(687,416){1}
wire [1:0] w11;    //: /sn:0 {0}(-27,-33)(-27,-23)(106,-23)(106,-10){1}
wire w2;    //: /sn:0 {0}(243,212)(204,212){1}
wire [31:0] R0;    //: {0}(77,228)(77,299)(41,299)(41,353){1}
wire [31:0] w5;    //: /sn:0 {0}(675,416)(675,372)(497,372)(497,228){1}
wire [31:0] w9;    //: /sn:0 {0}(663,416)(663,387)(309,387)(309,223){1}
//: enddecls

  //: joint g8 (w18) @(6, 122) /w:[ 7 -1 8 10 ]
  //: input g4 (Read2) @(-239,145) /sn:0 /w:[ 0 ]
  //: joint g44 (clr) @(353, -83) /w:[ 3 -1 4 10 ]
  //: input g3 (Write) @(-240,-38) /sn:0 /w:[ 0 ]
  //: joint g16 (clk) @(165, 285) /w:[ 5 6 8 -1 ]
  //: joint g47 (clr) @(541, -83) /w:[ 1 -1 2 12 ]
  //: input g17 (Read1) @(-239,96) /sn:0 /w:[ 0 ]
  //: joint g26 (w19) @(229, 106) /w:[ 5 -1 6 12 ]
  //: output g2 (Data2) @(668,482) /sn:0 /R:3 /w:[ 0 ]
  tran g23(.Z(w24), .I(Write[2:0]));   //: @(-65,-39) /sn:0 /R:1 /w:[ 9 1 2 ] /ss:1
  tran g30(.Z(w10), .I(Read2[4:3]));   //: @(-140,143) /sn:0 /R:1 /w:[ 0 1 2 ] /ss:1
  //: output g1 (Data1) @(59,462) /sn:0 /R:3 /w:[ 1 ]
  //: joint g39 (RegWrite) @(372, 263) /w:[ 6 8 5 -1 ]
  Regs8x32 g24 (.DIN(WriteData), .SD(w24), .SA(w19), .SB(w18), .RegWr(w31), .clk(w2), .clr(clr), .AOUT(R1), .BOUT(w9));   //: @(244, 153) /sz:(98, 69) /sn:0 /p:[ Ti0>11 Li0>13 Li1>13 Li2>13 Li3>0 Li4>0 Ri0>11 Bo0<0 Bo1<1 ]
  Regs8x32 g29 (.DIN(WriteData), .SD(w24), .SA(w19), .SB(w18), .RegWr(w4), .clk(w22), .clr(clr), .AOUT(R2), .BOUT(w5));   //: @(432, 158) /sz:(98, 69) /sn:0 /p:[ Ti0>13 Li0>0 Li1>0 Li2>0 Li3>1 Li4>1 Ri0>13 Bo0<1 Bo1<1 ]
  //: comment g51 /dolink:0 /link:"" @(395,229) /sn:0
  //: /line:"Regs 16-23"
  //: /end
  tran g18(.Z(w19), .I(Read1[2:0]));   //: @(-95,93) /sn:0 /R:1 /w:[ 9 3 4 ] /ss:1
  //: supply1 g10 (w21) @(68,-11) /sn:0 /w:[ 1 ]
  //: joint g25 (w18) @(210, 122) /w:[ 5 -1 6 12 ]
  //: comment g49 /dolink:0 /link:"" @(210,225) /sn:0
  //: /line:"Regs 8-15"
  //: /end
  //: comment g50 /dolink:0 /link:"" @(585,229) /sn:0
  //: /line:"Regs 24-31"
  //: /end
  Regs8x32 g6 (.DIN(WriteData), .SD(w24), .SA(w19), .SB(w18), .RegWr(w16), .clk(w1), .clr(clr), .AOUT(R0), .BOUT(w0));   //: @(40, 158) /sz:(98, 69) /sn:0 /p:[ Ti0>9 Li0>11 Li1>11 Li2>11 Li3>0 Li4>1 Ri0>9 Bo0<0 Bo1<1 ]
  //: joint g7 (w19) @(23, 106) /w:[ 7 -1 8 10 ]
  demux g9 (.I(w11), .E(w21), .Z0(w16), .Z1(w31), .Z2(w4), .Z3(w20));   //: @(106,3) /sn:0 /w:[ 1 0 1 1 0 0 ]
  and g35 (.I0(clk), .I1(RegWrite), .Z(w22));   //: @(394,217) /sn:0 /delay:" 1" /w:[ 3 9 0 ]
  tran g31(.Z(w6), .I(Read1[4:3]));   //: @(-123,93) /sn:0 /R:1 /w:[ 1 1 2 ] /ss:1
  tran g22(.Z(w18), .I(Read2[2:0]));   //: @(-93,142) /sn:0 /R:1 /w:[ 9 3 4 ] /ss:0
  and g36 (.I0(clk), .I1(RegWrite), .Z(w23));   //: @(567,217) /sn:0 /delay:" 1" /w:[ 0 7 0 ]
  //: joint g41 (w19) @(419, 107) /w:[ 2 -1 4 1 ]
  //: joint g45 (WriteData) @(479, 75) /w:[ 1 -1 2 12 ]
  and g33 (.I0(clk), .I1(RegWrite), .Z(w1));   //: @(-27,217) /sn:0 /delay:" 1" /w:[ 11 13 0 ]
  //: input g42 (clr) @(-237,-92) /sn:0 /w:[ 7 ]
  //: joint g40 (w18) @(402, 123) /w:[ 2 -1 4 1 ]
  //: input g12 (clk) @(-239,285) /sn:0 /w:[ 13 ]
  and g34 (.I0(clk), .I1(RegWrite), .Z(w2));   //: @(194,212) /sn:0 /delay:" 1" /w:[ 7 11 1 ]
  //: joint g28 (w24) @(381, 139) /w:[ 2 -1 4 1 ]
  Regs8x32 g46 (.DIN(WriteData), .SD(w24), .SA(w19), .SB(w18), .RegWr(w20), .clk(w23), .clr(clr), .AOUT(w3), .BOUT(R3));   //: @(622, 158) /sz:(98, 69) /sn:0 /p:[ Ti0>0 Li0>3 Li1>3 Li2>3 Li3>1 Li4>1 Ri0>0 Bo0<1 Bo1<0 ]
  //: joint g11 (w24) @(-15, 138) /w:[ 7 -1 8 10 ]
  mux g14 (.I0(R0), .I1(R1), .I2(R2), .I3(w3), .S(w6), .Z(Data1));   //: @(59,369) /sn:0 /w:[ 1 1 0 0 0 0 ] /ss:0 /do:0
  tran g5(.Z(w11), .I(Write[4:3]));   //: @(-27,-39) /sn:0 /R:1 /w:[ 0 3 4 ] /ss:1
  //: joint g19 (clk) @(-58, 285) /w:[ 9 10 12 -1 ]
  //: joint g21 (w24) @(193, 138) /w:[ 5 -1 6 12 ]
  //: input g32 (RegWrite) @(-239,263) /sn:0 /w:[ 0 ]
  //: joint g20 (WriteData) @(87, 75) /w:[ 5 -1 6 8 ]
  //: joint g38 (RegWrite) @(173, 263) /w:[ 4 10 3 -1 ]
  //: joint g15 (clk) @(362, 285) /w:[ 1 2 4 -1 ]
  //: joint g43 (clr) @(148, -83) /w:[ 5 -1 6 8 ]
  //: input g0 (WriteData) @(-239,73) /sn:0 /w:[ 7 ]
  //: joint g27 (WriteData) @(290, 75) /w:[ 3 -1 4 10 ]
  //: comment g48 /dolink:0 /link:"" @(11,228) /sn:0
  //: /line:"Regs 0-7"
  //: /end
  //: joint g37 (RegWrite) @(-69, 263) /w:[ 2 12 1 -1 ]
  mux g13 (.I0(w0), .I1(w9), .I2(w5), .I3(R3), .S(w10), .Z(Data2));   //: @(669,432) /sn:0 /w:[ 0 0 0 1 1 1 ] /ss:0 /do:0

endmodule

module Regs8x32(SB, SA, BOUT, AOUT, clk, clr, RegWr, SD, DIN);
//: interface  /sz:(98, 69) /bd:[ Ti0>DIN[31:0](47/98) Li0>clk(59/69) Li1>RegWr(47/69) Li2>SB[2:0](22/69) Li3>SA[2:0](11/69) Li4>SD[2:0](35/69) Ri0>clr(35/69) Bo0<BOUT[31:0](65/98) Bo1<AOUT[31:0](37/98) ]
input [31:0] DIN;    //: /sn:0 {0}(531,269)(531,318){1}
//: {2}(533,320)(627,320){3}
//: {4}(631,320)(715,320){5}
//: {6}(719,320)(807,320)(807,429){7}
//: {8}(717,322)(717,352){9}
//: {10}(629,322)(629,433){11}
//: {12}(529,320)(435,320){13}
//: {14}(431,320)(342,320){15}
//: {16}(338,320)(264,320){17}
//: {18}(260,320)(181,320)(181,352){19}
//: {20}(262,322)(262,439){21}
//: {22}(340,322)(340,351){23}
//: {24}(433,322)(433,436){25}
//: {26}(531,322)(531,348){27}
output [31:0] BOUT;    //: /sn:0 {0}(516,697)(516,672){1}
input [2:0] SD;    //: /sn:0 {0}(782,138)(852,138)(852,156){1}
supply1 w21;    //: /sn:0 {0}(828,169)(801,169)(801,153){1}
input [2:0] SB;    //: /sn:0 {0}(466,659)(493,659){1}
input RegWr;    //: /sn:0 {0}(48,363)(68,363)(68,378)(82,378){1}
input [2:0] SA;    //: /sn:0 {0}(256,657)(231,657){1}
input clr;    //: /sn:0 /dp:1 {0}(959,337)(1032,337){1}
input clk;    //: /sn:0 {0}(82,383)(68,383)(68,398)(55,398){1}
output [31:0] AOUT;    //: /sn:0 {0}(279,670)(279,702){1}
wire [31:0] w16;    //: /sn:0 {0}(531,369)(531,574)(520,574){1}
//: {2}(516,574)(282,574)(282,641){3}
//: {4}(518,576)(518,587)(519,587)(519,643){5}
wire w7;    //: /sn:0 {0}(472,451)(513,451)(513,405)(848,405)(848,185){1}
wire [31:0] R5;    //: {0}(288,641)(288,586)(525,586){1}
//: {2}(529,586)(629,586)(629,454){3}
//: {4}(527,588)(527,617)(525,617)(525,643){5}
wire w4;    //: /sn:0 {0}(943,337)(906,337){1}
//: {2}(902,337)(767,337){3}
//: {4}(763,337)(588,337){5}
//: {6}(584,337)(390,337){7}
//: {8}(386,337)(231,337)(231,357)(220,357){9}
//: {10}(388,339)(388,356)(379,356){11}
//: {12}(586,339)(586,353)(570,353){13}
//: {14}(765,339)(765,357)(756,357){15}
//: {16}(904,339)(904,417)(865,417){17}
//: {18}(861,417)(675,417){19}
//: {20}(671,417)(489,417){21}
//: {22}(485,417)(302,417)(302,444)(301,444){23}
//: {24}(487,419)(487,441)(472,441){25}
//: {26}(673,419)(673,438)(668,438){27}
//: {28}(863,419)(863,434)(846,434){29}
wire [31:0] R2;    //: {0}(262,641)(262,537){1}
//: {2}(264,535)(499,535)(499,643){3}
//: {4}(262,533)(262,460){5}
wire w0;    //: /sn:0 {0}(770,439)(764,439)(764,481)(579,481){1}
//: {2}(577,479)(577,443)(592,443){3}
//: {4}(575,481)(390,481){5}
//: {6}(388,479)(388,446)(396,446){7}
//: {8}(386,481)(214,481){9}
//: {10}(212,479)(212,449)(225,449){11}
//: {12}(210,481)(125,481)(125,383){13}
//: {14}(127,381)(291,381){15}
//: {16}(295,381)(477,381){17}
//: {18}(481,381)(660,381)(660,362)(680,362){19}
//: {20}(479,379)(479,358)(494,358){21}
//: {22}(293,379)(293,361)(303,361){23}
//: {24}(125,379)(125,362)(144,362){25}
//: {26}(123,381)(103,381){27}
wire w3;    //: /sn:0 {0}(835,185)(835,397)(330,397)(330,454)(301,454){1}
wire [31:0] R7;    //: {0}(807,450)(807,609)(541,609){1}
//: {2}(537,609)(302,609)(302,641){3}
//: {4}(539,611)(539,643){5}
wire w12;    //: /sn:0 {0}(756,367)(787,367)(787,258)(868,258)(868,185){1}
wire w10;    //: /sn:0 {0}(846,444)(875,444)(875,185){1}
wire [31:0] R4;    //: {0}(340,372)(340,545){1}
//: {2}(342,547)(505,547)(505,643){3}
//: {4}(338,547)(268,547)(268,641){5}
wire [31:0] R3;    //: {0}(512,643)(512,559)(435,559){1}
//: {2}(433,557)(433,457){3}
//: {4}(431,559)(275,559)(275,641){5}
wire w8;    //: /sn:0 {0}(220,367)(249,367)(249,213)(828,213)(828,185){1}
wire Z5;    //: /sn:0 {0}(861,185)(861,413)(700,413)(700,448)(668,448){1}
wire w14;    //: /sn:0 {0}(379,366)(414,366)(414,229)(841,229)(841,185){1}
wire [31:0] R0;    //: {0}(492,643)(492,523)(257,523){1}
//: {2}(253,523)(181,523)(181,373){3}
//: {4}(255,525)(255,641){5}
wire w15;    //: /sn:0 {0}(570,363)(608,363)(608,244)(855,244)(855,185){1}
wire [31:0] R10;    //: /sn:0 {0}(295,641)(295,600)(530,600){1}
//: {2}(534,600)(717,600)(717,373){3}
//: {4}(532,602)(532,643){5}
//: enddecls

  //: joint g8 (w16) @(518, 574) /w:[ 1 -1 2 4 ]
  //: input g4 (SB) @(464,659) /sn:0 /w:[ 0 ]
  //: input g3 (SA) @(229,657) /sn:0 /w:[ 1 ]
  //: joint g16 (R3) @(433, 559) /w:[ 1 2 4 -1 ]
  //: joint g17 (R4) @(340, 547) /w:[ 2 1 4 -1 ]
  //: joint g26 (DIN) @(340, 320) /w:[ 15 -1 16 22 ]
  register R5 (.Q(R5), .D(DIN), .EN(Z5), .CLR(w4), .CK(!w0));   //: @(629,443) /w:[ 3 11 1 27 3 ]
  //: output g2 (BOUT) @(516,694) /sn:0 /R:3 /w:[ 0 ]
  //: joint g23 (w4) @(765, 337) /w:[ 3 -1 4 14 ]
  //: joint g30 (w0) @(212, 481) /w:[ 9 10 12 -1 ]
  //: output g1 (AOUT) @(279,699) /sn:0 /R:3 /w:[ 1 ]
  //: joint g39 (DIN) @(262, 320) /w:[ 17 -1 18 20 ]
  //: joint g24 (DIN) @(531, 320) /w:[ 2 1 12 26 ]
  //: joint g29 (w0) @(388, 481) /w:[ 5 6 8 -1 ]
  register R2 (.Q(R4), .D(DIN), .EN(w14), .CLR(w4), .CK(!w0));   //: @(340,361) /w:[ 0 23 0 11 23 ]
  register R7 (.Q(R7), .D(DIN), .EN(w10), .CLR(w4), .CK(!w0));   //: @(807,439) /w:[ 0 7 0 29 0 ]
  //: joint g18 (R2) @(262, 535) /w:[ 2 4 -1 1 ]
  //: supply1 g10 (w21) @(812,153) /sn:0 /w:[ 1 ]
  not g25 (.I(clr), .Z(w4));   //: @(953,337) /sn:0 /R:2 /w:[ 0 0 ]
  //: joint g6 (R7) @(539, 609) /w:[ 1 -1 2 4 ]
  register R6 (.Q(R10), .D(DIN), .EN(w12), .CLR(w4), .CK(!w0));   //: @(717,362) /w:[ 3 9 0 15 19 ]
  //: joint g7 (R10) @(532, 600) /w:[ 2 -1 1 4 ]
  register R4 (.Q(w16), .D(DIN), .EN(w15), .CLR(w4), .CK(!w0));   //: @(531,358) /w:[ 0 27 0 13 21 ]
  demux g9 (.I(SD), .E(w21), .Z0(!w8), .Z1(!w3), .Z2(!w14), .Z3(!w7), .Z4(!w15), .Z5(!Z5), .Z6(!w12), .Z7(!w10));   //: @(852,169) /sn:0 /w:[ 1 0 1 0 1 1 1 0 1 1 ]
  and g35 (.I0(RegWr), .I1(clk), .Z(w0));   //: @(93,381) /sn:0 /delay:" 1" /w:[ 1 0 27 ]
  //: joint g31 (w4) @(863, 417) /w:[ 17 -1 18 28 ]
  //: joint g22 (w4) @(586, 337) /w:[ 5 -1 6 12 ]
  register R3 (.Q(R3), .D(DIN), .EN(w7), .CLR(w4), .CK(!w0));   //: @(433,446) /w:[ 3 25 0 25 7 ]
  register R1 (.Q(R2), .D(DIN), .EN(w3), .CLR(w4), .CK(!w0));   //: @(262,449) /w:[ 5 21 1 23 11 ]
  //: joint g36 (w4) @(904, 337) /w:[ 1 -1 2 16 ]
  //: joint g41 (DIN) @(717, 320) /w:[ 6 -1 5 8 ]
  //: joint g33 (w4) @(673, 417) /w:[ 19 -1 20 26 ]
  //: joint g42 (DIN) @(629, 320) /w:[ 4 -1 3 10 ]
  //: joint g40 (DIN) @(433, 320) /w:[ 13 -1 14 24 ]
  //: joint g12 (w0) @(479, 381) /w:[ 18 20 17 -1 ]
  //: input g34 (clk) @(53,398) /sn:0 /w:[ 1 ]
  //: input g28 (clr) @(1034,337) /sn:0 /R:2 /w:[ 1 ]
  //: joint g11 (w0) @(293, 381) /w:[ 16 22 15 -1 ]
  //: input g5 (RegWr) @(46,363) /sn:0 /w:[ 0 ]
  mux g14 (.I0(R0), .I1(R2), .I2(R4), .I3(R3), .I4(w16), .I5(R5), .I6(R10), .I7(R7), .S(SA), .Z(AOUT));   //: @(279,657) /sn:0 /w:[ 5 0 5 5 3 0 0 3 0 0 ] /ss:0 /do:0
  //: joint g19 (R0) @(255, 523) /w:[ 1 -1 2 4 ]
  //: joint g21 (w4) @(388, 337) /w:[ 7 -1 8 10 ]
  //: joint g32 (w4) @(487, 417) /w:[ 21 -1 22 24 ]
  //: input g20 (SD) @(780,138) /sn:0 /w:[ 0 ]
  register R0 (.Q(R0), .D(DIN), .EN(w8), .CLR(w4), .CK(!w0));   //: @(181,362) /w:[ 3 19 0 9 25 ]
  //: joint g38 (w0) @(577, 481) /w:[ 1 2 4 -1 ]
  //: joint g15 (R5) @(527, 586) /w:[ 2 -1 1 4 ]
  //: input g0 (DIN) @(531,267) /sn:0 /R:3 /w:[ 0 ]
  //: joint g27 (w0) @(125, 381) /w:[ 14 24 26 13 ]
  mux g13 (.I0(R0), .I1(R2), .I2(R4), .I3(R3), .I4(w16), .I5(R5), .I6(R10), .I7(R7), .S(SB), .Z(BOUT));   //: @(516,659) /sn:0 /w:[ 0 3 3 0 5 5 5 5 1 1 ] /ss:0 /do:0

endmodule

module FETCH(clk, PCNew, Reset, Inst, PCNext);
//: interface  /sz:(113, 114) /bd:[ Li0>Reset(33/114) Li1>PCNew[31:0](66/114) Li2>clk(96/114) Ro0<PCNext[31:0](36/114) Ro1<Inst[31:0](88/114) ]
supply0 w6;    //: /sn:0 {0}(571,436)(571,414){1}
supply0 w4;    //: /sn:0 {0}(472,348)(472,329)(454,329)(454,351){1}
input [31:0] PCNew;    //: /sn:0 {0}(383,389)(438,389){1}
output [31:0] Inst;    //: /sn:0 /dp:1 {0}(686,387)(588,387){1}
output [31:0] PCNext;    //: /sn:0 /dp:1 {0}(689,299)(623,299){1}
input Reset;    //: /sn:0 {0}(381,328)(444,328)(444,351){1}
input clk;    //: /sn:0 {0}(404,455)(449,455)(449,427){1}
supply0 w5;    //: /sn:0 {0}(574,254)(574,244)(608,244)(608,275){1}
wire w13;    //: /sn:0 {0}(608,323)(608,338)(625,338){1}
wire [31:0] w0;    //: /sn:0 {0}(475,256)(475,315)(594,315){1}
wire [31:0] w1;    //: /sn:0 /dp:1 {0}(553,389)(516,389){1}
//: {2}(514,387)(514,283)(594,283){3}
//: {4}(512,389)(459,389){5}
//: enddecls

  //: supply0 g8 (w4) @(472,354) /sn:0 /w:[ 0 ]
  rom g4 (.A(w1), .D(Inst), .OE(w6));   //: @(571,388) /sn:0 /w:[ 0 1 1 ] /mem:"/home/omiralles03/Documents/Estructura de Computadors/Practica2_EstructuraComputadors/TAREAS/mult.mem"
  //: input g3 (clk) @(402,455) /sn:0 /w:[ 0 ]
  //: input g2 (PCNew) @(381,389) /sn:0 /w:[ 0 ]
  //: input g1 (Reset) @(379,328) /sn:0 /w:[ 0 ]
  led g10 (.I(w13));   //: @(632,338) /sn:0 /R:3 /w:[ 1 ] /type:0
  add g6 (.A(w0), .B(w1), .S(PCNext), .CI(w5), .CO(w13));   //: @(610,299) /sn:0 /R:1 /w:[ 1 3 1 1 0 ]
  //: supply0 g9 (w5) @(574,260) /sn:0 /w:[ 0 ]
  //: joint g7 (w1) @(514, 389) /w:[ 1 2 4 -1 ]
  //: output g12 (Inst) @(683,387) /sn:0 /w:[ 0 ]
  //: supply0 g11 (w6) @(571,442) /sn:0 /w:[ 0 ]
  register g5 (.Q(w1), .D(PCNew), .EN(w4), .CLR(Reset), .CK(!clk));   //: @(449,389) /sn:0 /R:1 /w:[ 5 1 1 1 1 ]
  //: dip g0 (w0) @(475,246) /sn:0 /w:[ 0 ] /st:1
  //: output g13 (PCNext) @(686,299) /sn:0 /w:[ 0 ]

endmodule

module main;    //: root_module
wire w6;    //: /sn:0 /dp:1 {0}(778,326)(778,341)(750,341){1}
wire [4:0] w13;    //: /sn:0 {0}(229,345)(152,345){1}
wire [31:0] w7;    //: /sn:0 {0}(823,436)(441,436)(441,381){1}
//: {2}(443,379)(497,379){3}
//: {4}(439,379)(404,379){5}
wire w34;    //: /sn:0 {0}(22442,-11681)(22442,-11671){1}
wire [31:0] w39;    //: /sn:0 /dp:1 {0}(526,389)(588,389){1}
wire [31:0] w25;    //: /sn:0 {0}(750,379)(782,379){1}
//: {2}(786,379)(823,379){3}
//: {4}(784,381)(784,494)(969,494)(969,412)(1013,412){5}
wire [31:0] w4;    //: /sn:0 {0}(83,327)(146,327){1}
//: {2}(148,325)(148,309){3}
//: {4}(148,308)(148,268){5}
//: {6}(148,267)(148,145){7}
//: {8}(148,144)(148,140){9}
//: {10}(148,329)(148,344){11}
//: {12}(148,345)(148,443){13}
//: {14}(148,444)(148,461){15}
wire w0;    //: /sn:0 {0}(688,90)(734,90)(734,117){1}
wire [31:0] w3;    //: /sn:0 {0}(83,275)(118,275)(118,175)(670,175){1}
wire [31:0] w20;    //: /sn:0 /dp:1 {0}(1013,392)(955,392){1}
wire w29;    //: /sn:0 {0}(22476,-11710)(22476,-11700){1}
wire [31:0] w19;    //: /sn:0 {0}(404,447)(464,447)(464,401){1}
//: {2}(466,399)(497,399){3}
//: {4}(464,397)(464,209)(670,209){5}
wire w18;    //: /sn:0 {0}(349,478)(349,508)(-65,508)(-65,274){1}
//: {2}(-63,272)(-32,272){3}
//: {4}(-67,272)(-77,272){5}
wire [4:0] w12;    //: /sn:0 {0}(229,309)(152,309){1}
wire [31:0] w23;    //: /sn:0 {0}(588,344)(404,344){1}
wire w10;    //: /sn:0 {0}(315,238)(315,228){1}
wire [31:0] w24;    //: /sn:0 /dp:1 {0}(1042,402)(1066,402)(1066,556)(197,556)(197,413)(229,413){1}
wire w1;    //: /sn:0 {0}(523,316)(513,316)(513,366){1}
wire w31;    //: /sn:0 {0}(4281,420)(4271,420){1}
wire w8;    //: /sn:0 {0}(747,252)(761,252)(761,225){1}
wire w27;    //: /sn:0 {0}(1016,456)(1029,456)(1029,425){1}
wire [31:0] w35;    //: /sn:0 {0}(790,170)(831,170)(831,64)(-52,64)(-52,305)(-32,305){1}
wire [25:0] w28;    //: /sn:0 {0}(670,145)(152,145){1}
wire [3:0] w14;    //: /sn:0 {0}(641,260)(641,292){1}
wire [4:0] w11;    //: /sn:0 {0}(229,268)(152,268){1}
wire w2;    //: /sn:0 {0}(-32,335)(-52,335)(-52,547){1}
//: {2}(-50,549)(287,549)(287,478){3}
//: {4}(-54,549)(-85,549){5}
wire [15:0] w15;    //: /sn:0 {0}(229,444)(152,444){1}
wire w5;    //: /sn:0 {0}(880,347)(880,337){1}
wire w9;    //: /sn:0 {0}(867,522)(888,522)(888,473){1}
wire w40;    //: /sn:0 {0}(190,379)(229,379){1}
//: enddecls

  //: switch g8 (w0) @(671,90) /sn:0 /w:[ 0 ] /st:0
  JUMP g4 (.Jump(w0), .SignExtOut(w19), .PCNext(w3), .lnm26(w28), .PCSrc(w8), .PCin(w35));   //: @(671, 118) /sz:(118, 106) /sn:0 /p:[ Ti0>1 Li0>5 Li1>1 Li2>0 Bi0>1 Ro0<0 ]
  //: switch g16 (w1) @(541,316) /sn:0 /R:2 /w:[ 0 ] /st:0
  EXE g3 (.ALU_OP(w14), .B(w39), .A(w23), .Zero(w6), .Result(w25));   //: @(589, 293) /sz:(160, 125) /sn:0 /p:[ Ti0>1 Li0>1 Li1>0 Ro0<1 Ro1<0 ]
  //: joint g26 (w18) @(-65, 272) /w:[ 2 -1 4 1 ]
  //: joint g17 (w7) @(441, 379) /w:[ 2 -1 4 1 ]
  READ g2 (.RegWrite(w10), .RegDst(w40), .SignExtIn(w15), .WriteData(w24), .Write(w13), .Read2(w12), .Read1(w11), .clr(w18), .clk(w2), .Data1(w23), .Data2(w7), .SignExtOut(w19));   //: @(230, 239) /sz:(173, 238) /sn:0 /p:[ Ti0>0 Li0>1 Li1>0 Li2>1 Li3>0 Li4>0 Li5>0 Bi0>0 Bi1>3 Ro0<1 Ro1<5 Ro2<0 ]
  led g23 (.I(w6));   //: @(778,319) /sn:0 /w:[ 0 ] /type:3
  //: switch g24 (w8) @(730,252) /sn:0 /w:[ 0 ] /st:0
  MEM g1 (.MemWrite(w5), .WriteData(w7), .Address(w25), .MemRead(w9), .ReadData(w20));   //: @(824, 348) /sz:(130, 124) /sn:0 /p:[ Ti0>0 Li0>0 Li1>3 Bi0>1 Ro0<1 ]
  //: switch g18 (w31) @(4299,420) /sn:0 /R:2 /w:[ 0 ] /st:0
  //: dip g25 (w14) @(641,250) /sn:0 /w:[ 0 ] /st:0
  tran g10(.Z(w11), .I(w4[25:21]));   //: @(146,268) /sn:0 /R:2 /w:[ 1 5 6 ] /ss:1
  //: switch g6 (w40) @(173,379) /sn:0 /w:[ 0 ] /st:0
  tran g9(.Z(w28), .I(w4[25:0]));   //: @(146,145) /sn:0 /R:2 /w:[ 1 7 8 ] /ss:1
  //: switch g7 (w18) @(-94,272) /sn:0 /w:[ 5 ] /st:0
  //: joint g22 (w25) @(784, 379) /w:[ 2 -1 1 4 ]
  //: switch g31 (w29) @(22476,-11723) /sn:0 /R:3 /w:[ 0 ] /st:0
  tran g12(.Z(w15), .I(w4[15:0]));   //: @(146,444) /sn:0 /R:2 /w:[ 1 14 13 ] /ss:1
  //: joint g28 (w2) @(-52, 549) /w:[ 2 1 4 -1 ]
  //: joint g14 (w4) @(148, 327) /w:[ -1 2 1 10 ]
  tran g11(.Z(w12), .I(w4[20:16]));   //: @(146,309) /sn:0 /R:2 /w:[ 1 3 4 ] /ss:1
  mux g5 (.I0(w19), .I1(w7), .S(w1), .Z(w39));   //: @(513,389) /sn:0 /R:1 /w:[ 3 3 1 0 ] /ss:1 /do:0
  //: switch g21 (w9) @(850,522) /sn:0 /w:[ 0 ] /st:0
  mux g19 (.I0(w25), .I1(w20), .S(w27), .Z(w24));   //: @(1029,402) /sn:0 /R:1 /w:[ 5 0 1 0 ] /ss:0 /do:0
  //: switch g20 (w27) @(999,456) /sn:0 /w:[ 0 ] /st:0
  //: switch g32 (w34) @(22442,-11694) /sn:0 /R:3 /w:[ 0 ] /st:0
  //: joint g15 (w19) @(464, 399) /w:[ 2 4 -1 1 ]
  FETCH g0 (.clk(w2), .PCNew(w35), .Reset(w18), .Inst(w4), .PCNext(w3));   //: @(-31, 239) /sz:(113, 114) /sn:0 /p:[ Li0>0 Li1>1 Li2>3 Ro0<0 Ro1<0 ]
  clock g27 (.Z(w2));   //: @(-98,549) /sn:0 /w:[ 5 ] /omega:100 /phi:0 /duty:50
  tran g13(.Z(w13), .I(w4[15:11]));   //: @(146,345) /sn:0 /R:2 /w:[ 1 12 11 ] /ss:1

endmodule
